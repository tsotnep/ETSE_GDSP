library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use work.txt_util.all;
USE ieee.numeric_std.ALL;
use work.MATRIX_MUL_IP_CORE_LIBRARY_Syn.all;

package MATRIX_MUL_IP_CORE_LIBRARY_Sim is




-- procedure print_memarray_data_output(Data_input: inout std_logic_vector(DATA_WIDTH-1 downto 0); clk_period: inout time; stop_signal: inout std_logic);
-- procedure PrintResultToConsole;
-- procedure PrintResultInCSVFormat;

end package MATRIX_MUL_IP_CORE_LIBRARY_Sim;

package body MATRIX_MUL_IP_CORE_LIBRARY_Sim is


end package body MATRIX_MUL_IP_CORE_LIBRARY_Sim;
