XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5��x^�p��i�;�78�"f��@t���������ʜ��Y�p*{S����e�x�]�T�%[G��e���3���򔽩9���u��ehz_I״�l��Zbq���o��Gd��yaC�T�`���ϔ�>�������`5�T�%c�<8�6�,� ��ОIɸ�(�@F�Mo�1��ѿ�x	۟5��7���U�ˌ����P Q����^������ɦ���N�V��iٳ�Q�A��l��# �FE��?I�W�<v9im���"�r��� _!(��7���L���p����<�K�p�<�Zߐ�yj4
����5�{�XA��n\��Z�
�(�7e�M�����������?�H��,Qr�"��dɎ�UUڰg�M� a��i�B���q��9��f���m�����W~�u����Ń�w��Z��[P�"�$��1��&��_�	W��FDg�`�&3kS��>�B%8����Y�X4���R��ʨ��?�DZ�qò�>@SRD�'Q������a���G ��0��uA��4ĥhs�OJ&)�rn���Ͷ�4a;�����9�N���\`Zy	��FkSǋ�IGf(�y����z���z�j/�k�C��\�u�Q���ίI����[X���2�n�D�� �k���w����NT�_�|�
�UK������}Λ2�Yh#OS{<:� 8^�]��dGosB�s�oͪQ��J\��5�ZΏ���ܴ�t�/b���^�XlxVHYEB    aa52    13d0�2r��`��y��>u���Fb��0�Vj�9�i��w\�l�v'fL�C�b�f�	�5>�c�)�����.�-�W�Sh����p��} 8�����+��%iX Yĕؗ
!���fpX�6���G����_ٹ��~7	��}��"Hr����
�p[ON�l*�:]R%I(�d��'�����y"Lb�&��u�ʈ���o*>kƞ�Ű&wx�g��1e���w<7�������ڙ����ؗ��z�V4T}�n��
���(ґ@��_����3��#_��^��);Эx�V����[M�۶v-�ٛ{����E��t�Kq���4�؇�-w�G�������P�4PBJ.Kө��c���c=$b��̧�6؆�����.v�3sk�p����`k>����y���B^Npø�$��V�[4C��tP@�ͼ��C�:[�!����yg,*#Ok�ך���6t�v�X�����
�]f�k���U�rw�Vw��p�;���4O���F~��B䣂o豲��js�<��"�É��l8�p!ī� ���\��{��]�=z���F���/G�I�jx�"U1��ʈ���P+P�����r6���I��u��8��B����+F���J9�I.F�H|P��,�	n9aC��f��E����O�X�?u3�^�x?ܬ�cf��̀ p�f���|Zф�q�T:S2�H lo����<��q[��<���R4_qC��yQF���[���?�8ʚ
Է�9dF6��m��?��/���(�g�brs�wJ��ݏ;틕��\����6C�1��x3�3�n>O�I�������?�u���Rn7�2}�$�Kg�j�VZ<� J�D� m�nu) �i@}@rgʶ�E�O9j�c^�qq_�M�Y���S�E���.�q������xy��>�]��?�ŗ2�)���Vd��� ([�IJ8oI[�������yA�iH����CO�K)����z��4� �|7d�ܥ����Օۡ��c�.H|��t%���]J��1�UqҒ���n�U�� ��@�)���̩��?XV���Z+L�425~j �D31�X���u��U��h���ט�Xܮ�TQ�%�g�K�Ɔ�O�|����&��P�!�U�Յ���*���=J��j^�xڡ�K����>5�f�����]��BG�9T�{��:0pey�Se�%
��>�n�\M���J��ׇ�P� �]��΁���ߧ� �Y���zc���/U�aX3 ��Ia,reI���o�2|�8���P*���q�ʽ��3�d���T&o��[�E�N�B���:�������5ѭ2IbY�y��Cl!�̝��N��I���|S2�d6~����y�+
M���9q���h�M��5�Z�v���0��,6$� �GW@o��*���Pbh�ɳ��6��Y�A�"��h O�F��ТM糶ݲ@"J#��~T�=�{\I�T�;����{�� ��K�o��^j�@�����[��"�#a�	�
s�h�xwJa�[=�������Y�K�r�7��M��l���f8i3< �?��1�zk�G���b̷]��qcX=�
�?�w�:pƏ�\N$�@�t�s��l�OΨoC��	.�LМ�IEM1IӺd(��z@j��pd��H���)�+6	��a�	ߎ�Go����mUՐנW����,�L�E��A���>x�e�%
��կ�`�:��I����O�P*�,})���������m^���C�C-	p͔9��������X��{n]gU��Vh�w��Rf	��-�cfV�M�m��]\��-�����}����sp�pJ}]01�X�D����˜���>g9v1�^���%�������J�.~�Df`ɬ�O<���U�N����[g3S�1]�?J#$NX�=p�JǯwV�2M�a��/��7#�o&��^��Y�x%�U��蜙�������2���鮺�9�_؞��+Y�K8QFn<�F����݌ΞyI�a�F�ݦ� C�fd���+�ECM���1�x� 	6�.�gy.��0�ȌtAƐIS.q��-���Dx�6V��.SAQ��J H��RHa���Q�U(�Ѷ� �M[����Ea}�#.1�������mt�m�]�77���)���v'>�`?N-��1R��e\���/�����/�F_+fH ������y��n�?8	[��"����I����%NK=ת.����3'�Vr��څ"\�l�-;�
�5�2|KW��Q�|H5��Am���q�^̔p��e�u�(_ke.8m��s�'����P������C��߉��p~A���V���KD�o���E&y��W[nŐoLNgLR�͏H$�aT��\R�t���$)���-HN�l;�r�I�s�Y�M�2���Y�Yw�$k�f8��{0���ko,�_8�tb�]Ȩ4`���G ��CZV����O��S�f��]~�+U���5���2!B��z7��sI	}��vH�
��b}Y2 D�pQlF<�+5�vN?��f ߄0�n>�Ç�;��JR���Dzu�󸲰�^��Z�t6��.ڤR���2�7֧�N�������K {�⨬��Bl�,n�b�^��>�X�dǃ&�9��?��Mb��0l�8�d���zDyY7?��DC��q�E��ś��~��L�:��(��`����i]=��5-��{'�2���>2��:��81�U%���ї_F}Яn)�W�n��1�욘v�y�d��-Rk��(���Z� ��.JɕY�b�t�-@[�t�����>�}�I��-#��T�5�Q׺r�4��KZ��&�)�����%X��o�,��3DOi,�h�����w�Gү��D$���m��\㥤��?�>�������	ò����<j�#�� J'ʅ
��4'����	>"�n��M�X�镞h�)�ڪt�MLQ!+H��Mv��]�d@#�u���M��d<� -n�IC��.��4�Ώ�c(�\"L�y�6F/ZD����jL&�!P����u���+��qȳ��议�+� t�ym�f���t=I��W*L΢��u�w8���[/�ɟ�0%��֖f*��⾞��1���{$�雯���li���Y��D��Ua��6�ѕ0��j��"m^�c���:�@ңd!�2�r������ρR��e'q�/�����Ä͉�c�)�M��
�i�ZZG�HT���Q��鲧7a�$>��r~�)��l�(mF��* �v�r��z���e�T4m�]ޒ��	�ӣµ�(�^]�QՑ��4�/q#��	�!3i��x��g�Ik쐐o ��M;	?���T[_��r�b�i�]�QS/˜�������iDy<a����,����K�6�_E��")+���;���oxz��Wy \l��:w:��")Be�Y�E\�]���fe"|�ַ��mDF[22���#����=�ٜ<Ea�%#�c--1e7��a���Hol�TWF_JR������J �`�<��L&�֠��J$q����{��6�� �yi1�ۋ��d�4�������&��'�(J��\#R�X����*X2Ym5�Ԏ��&),����'dϹ�M�R؆���M4!���5���8"hm���l׫Մ�)K@��JP1F
��޼͸fs�9HI�(�>�HCy�ɕ�H ����˫SA:x�y{�%!k�Xd$&\�'�!�$���-=&h����ДǤKy6���!�=�]���i>I����葚�te�ޤǵGw����Wɋ�xR�����B�ϳq�)�&	�"��ݤS���p��
S.�Î!7����,��5�g���|�C�}~U����drw:�yO/ɀq|eTX'Z���ԱTc�m��'�K��ɲ]��ͭ`�.k�2p �o]1�QO��a���˱�&��x�T=o,�?�h8�c����)�~����,�!tc�`�������./s�� ^m�=hr!�@��Y���b�l8�K)I����#��A��&���v�P����R-�m�����!� �8�~��Hք��+��Y�"�m�>�`a`W)�O��wƷ2�m�0��@bv�ˏڮ�+�t��w�֖�!�0l�k��e�N&�~�?�r��6�snbh���M�<�j��+�P#�� �����[M3�d��Oy�u�wC��H�,v��c��R:�N�uP��r ݩj��m0��n<�{Tf�#:���Q�B0�W�/�p]1���I�E��B�cX��?�K�t/m�=�b�rr*W���L�_1٤���Oѐ"K0-t���2��v�7�?0U����lV�8H��1�O��^���%�����r ��p櫔iմ g?bI�ط�!�]�o*��FY�9X(���ֺ���e�`�ܡ5�̲6�J�5_��d��ੵ��m8 ݐ�"��*ĺ�x��̏ɯ�9f����-TȆ�g����0�����������OO��1v�	����wp5�����@��s����.���4���G&=̙���P~
��Z�h+����@>Z>�F�YR�µ�����{��6ꌠ�'!���|
�X	��4�2��D���L���M�?�*Q/#ql,S�`��@�T�D�+T��[���1��h-�Z�,��U�r-4��
ر/��U8?��'�G�_;���qa�IîPjĎ ��g����^^Z'��<�����������;��rʃu��h��<a�i�;+f�V$��R�n�̙�m��I�걜V�t�^/<xr�l���T0`������@�s>��iO�E,��w_�S���?o�B(�EF%�cQR�����ב?b�U�� �H���US�-�&t�(���}��c���y�1�p�+�F�����J�FʙH�b�o~P1nSb�i��Wj���rmO��"�%I�9��D�63�B��6�b7��E�c�AC��e��Q�ET�7���-�*f�