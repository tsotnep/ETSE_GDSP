XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�býܤ����|S����P�2�Pw|��G�/�qv���703k�>�/�,��yL�K�#�����h�I�:��^��k
l叁Xi��L�����p;�O���_�A��1��O�������	=��	� g$Lv�6��5�><U&2�=�������vI��Cb/��6e���o(2�
�u�˕�d��K�XC�<���|~����Y�
e����<��1�?���E��eD��]�����9;f��6ҡ���7����nÃ�ߣ�*<h��;��{Ty�5e������o'Xb�`�'D���Q��G'�(xN4Wq׹�T�$������;��#?[{�iX$U3w){T�q-���.��-S�09A#0B{, �K��6.�(b�b���]%� {���_ɟ��VS!_P����@�IߖC)4!.�q���=�G�+�8��0�2@j>�s�`x��־JsJ÷iI�j�Tmj$�$���2�(�/&���%Q����o�_8�3|G�5�*9i��ߖ��O��#����F�Pd�y��X��!p
t�V>F��Z��#�i��ϷXoc���(3gٔ脮Th��#��52�ֿ��v$AYx�m�B'�P�gRD���S�_H_4Gi�!b���aX��R<}S*S�L�Q�t�[�6.sH�S8�������B�ɿ�4iވQo_���1�IV�	r�E,�;���<_>œ�:�F#tBr��RhO����!@�h�1�7a���7A������1�k�������(XlxVHYEB    56d2    12a0��r)�0��e�&��jÇ͍�a�1x,�WV5}Y/-b�Qԥ �sY~�B�tg'�KE�:��H�+�pi/��aΉ��>o��Ǝ�0^0�j��Ӌ�Q<�|3-t#����a�A�鉪����5�E;X�q��)}6Tf���rMCꢥ�%1̳1@�Tg1�'t�p�	�H���=oM>o���o(u�g��m�Ze�C��eݤG&%�Sħ���R�[Dc��eae�Pp�����o����xf� �8�"�v�U������c� a�����5���M�hG[&ʴ���6)E���+ӱ�Գq��eF�Ӏs� >�,�1�	���V��2F���sf���Q>������v_x�\����	�V�c�}5O�Yfv��v�8��;�+���ˣ�=0�]��G��x �z�;��́ct�
���ڽ&�$��r8�[-a% &5{7z�'c0焪0�V���-I}��N����oZ�f�rV��j��6�o �/@!��"(�>��$��+��P7;�|u>� ��u?Aq�|�R�����d��A7��Sxɗ�ͥ�p�)��7~�D(f`y��ǖ� ĵ�H8lUe�o� �]��;Mظ|�k��*��:�#H�
��.��q�|�<�K#�|zf�'��Ӡ��H_�_�:�Nc���ũ�G�,�HbF�vB1j���W�<�ӀIB¤s��O�;�`�,����;�3Y
�dgR������TX�� <0��HLX���ێ�K��E�8Fї��W�8z{(N����N|X5�`�\�*I���V/j!� ��X���}���gx�@8N�"*�*�&���I�E�(�h���B���,?�B���IޥǾ�����_��Y�V��S�ZM�b�\��Gs:c�����#���Nv5�@��f��k�z$��Y�VA��oͫ��khɘ��k]��$	:zZ1���m��(���w�s�:(5��+lMRc�)�3��ȯ���Z.��g��O_�Ti0`�AR�̝%R\<'��74��"I��eh:� S��}��r��j�"yc��c2F�B�ȏ��e�׵�#�ϳ��/
Zg�	�D�n�P,Kjؘ��\�D��B�B��9�'�D����K��\A�_=;|mzo�.�q�}�~H���wAQҥ3|��R��)8��az���wu��>a�(�v���D���ֆ�wb�g�N��g0e[$9~���C*n�V�q��|����
J�������k����/�<&5�)*۹�2$�.Ћ���N�Z7oc��̯�[֛zq����
C�J�۫S�����N(�SH�2���=`�@?U���H�7���k�3��t�/��2oT�@��z�;���Î��Ǿ�<�?e[�X�$*]��u�Y�En1z��}�v=���nȯ�л0仄��=�5A��&���{l��L�Ĥ|W��i N��K	��P)���Ye}>���;���9��(�Z�ƥ:�'��E�#��f]}��\�A��ϻ4�\�9�&�"Ɍ'S0��h�Tt!,H�)/�s�r�J�G��?-<I�'�q�t< �#L*���0J(�}�r�F�3�;F�(HJ��������n^��G�#��Y|������$(I�E��)��`�~�X<��y���B�v��N.զh?C߁���gp*�Ic4���^kk<�:@��uP���r,d>D��֮�,�f ��j�ѩ�* \syB���L"����Ϳ)D���<��Xc�5ˣ'�uJ��_�H�T#Wf�\	�n46�z>z�h��q%��1/����!
A�:���u�A�$X��� �V�x)v��*#Lk/�ٳܳͧ�>�C"�&�,�H�l���zr � z�􂷳�9ٿq��Lb�D�*��i\�e��L�H&A�{%����}'���5
ۓhr`�[ѷ!�a�����&"�[K)��wL�H!,R�_������/����j7ε���Ah�{�V!E����d��uDP�x�Vh(h�	�95���r��PA��/�G�YG�X��z���}��;��kйU�M�T�p-�v�ٵj���L2 ?����P���2�M�ňI���=#��S!���`�m���K|U��W^�B˳����l�
|���X[�X��I}���=vf��?W���i&�)�! N;"�G��}�F_'�99��*�R���~�ŭh	���œmzHpܱR9X�~�Cfo�^�d%�����J⺎�辗~���\��.-<����R5�P����h��뗔:fP_ Zn��q�<	�h���c��`|u)��ɈDx�����n�SwZ����yQ1��9+�qZY@�=�D�@�5�l�d���a�O,K�π�b]S~,J��z�e���?�i�M���K�0,iS��4��_�c!ƈ��Z���_�;�lϹw+�:΢���)��d�]%���"�i5�Чd�Ji���vFlm����5ح}]�<�dy{7fy OsV�����OA�(�r��Κb�w��8o*-s2n�;��?��|��Un]�7�wj�J���G�n����H�F�g�����)�dU-�d
mX=�	f<}T�C��fT�l\𕭚L3�>Y�`��Ҭ7�,�R�za���A�(��<����;&�ة.���Q��9+b)�t1&y�V����м���WC*�E&�ڋ�&^2]��ݮ����00���d+KJ|B)G��'�G���`6 [�9.k����H1�91J;_�qp�sx��w��U�Nf���?P��`�8�+�Le�qXk6KD�1.\B�ý�$v��\錘WE��X7�_��=��Lg���u*��;e,��&�[�R�<������V�X��j�`3g����<O��f�,�Q�5H+{f��Eb�?<c���r<Y��ݞ�v��FL�0HN�����F��j&��H�Q�D������]tH#|R�%�<L�:TU�l����U���A�/����a���`�H��%��M�J�7k1�U�.��c_oU@jܹF�Z�^��?�;;��$>��2��:����i�.�Ђe��YRk�Ơf��ߩ ��c�QE'ŬW��������͍w T)=G|)Z����7 #�ܡV��$Z�A� @)&����GJ?�A�08�;��/2�8P�U��v�x9�Ȇ��x���\Q�R���$��a������$�&��oP ��)i������|�N|�^�$iIA��+��3]>�a����{�ٹ�8��!h*r˔g���]v�E�.Ay��Hy���D�氇��s6b'�ZM<}�}+�h��Y]�)��3s�rt�m�����M⪬FUm?0��k��|hQ�����^j��i�[�p�.�"
0�^�etʳHW^M���5��2�? �8��>>�Sr�>~�������Ǉ��
��v���>�I\��x̏�Ѹ����p�����ϋT��|N>�$��B�DJ"Nj�l+-�N��c[ְ�lŭ��Y�a�T(=u�>�j�l��ƽ#�vM}�Gߏ��&S��E!2�f__�m ������1�Ç�See�)l��Lm��,v���S���$=���1�ey��퍕�H\*��Z��(Ru����k��e�k��,Au�C�Ӽ�݋����	&�b1z2���0�3m��H�ȵtn�k\~��,��l���� e���l3v.�f}�뾌"�����!�C3�'�P>�r�3�Z�##BB֧�G��'���ڠF�kL�\��Lqk�T`C����Z�q��~�e_ _�_H_[�h�5�:��3Pm-��@aW���e �[�Χڒ�R���}  �% ���$}�~��6���<jl���J?�v� �t�d[�ǻ�xX5+-34s�S�Z�X�_A0��C�ժ�|0حl#,�|�_�<e�_�!�7���e8�t��,��t_<=��	(
�B��>Vq&�A���I�E��J��+�7��ޒ�̾�T,�qU��HJ�b ��`��{�blb ���`���������J9�s0W�?�\��&)�#o�
��y�վd�Q�sզD�O�3㼓^�/�����	�in�W���J�4)�YM������JS}�v'�ք|c���tH޹B����$Ѱק$�\ՐP	֡���������[����26ѦOǗ���Q���D�S<�F�&�ot�$Q�n�j˯�,%R�5w�D9�+���դ����gv��>|B��_�Y�v�Q�L�gFt�ycQ��,L_3$QRț�e���}��I���:3���pH�$���6�^H GHv3��ǰLW�Rq��^�`�%��f��%+�Q��_
�{KYؠ,H��R�hrc�Z�kW@ ק�?�,�1S��d���/\��s�d��X�O��8��<Y��L3���g���GJ���o��8�թ��Kű0�mVy-��|8u���O�l��?�1�~��/��rMw�����<M����HN���FOHb��Iܦ&�$a�7K�a���o�D�OLI�8����hj���'������Q�UK����/స�-Q�Ӕb��4�,���Bń��"� ��F;f��8G�=oK����%�C}����p}�I�I8.u��i�;6�ܯgi�4�m��@u�-uNFϚ!穷���|z�nO�)���'#`W:�f�0���oSR�O`k��^�H`���F{u��6-�r���	C�M�����ƾ���'!�P*]�<\�~�0�"�Y�lu���r�;�$N��