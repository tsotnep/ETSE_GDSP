XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Sl^]���v7î�[��/`�eHs`县�wa��ķ]�홟�^f�B���^ �;;�O��,{I�9�m8D(�{�f�.#?Tή/�_)ދ�~��a�ZH���<�:�*6�EdΒ�'�fq.���7p
�cx��?6q����w+jA� B3��H~�a����+H�aG=�������]��Y|	�*=dPJE[-bZ�X&>8U%�;kt�zF���I?��!'5ݫo�@͹�c�l��Ċ��U�!�5��Bm���bp-�n����AN�O���5`'#�̤��h�/��~�t��(��I�����s�U]}��sV.��Y앐��>-�@[�m����r���FG��*@WP&r$��0ef?�l0���/˥�gU�m�ngS}>P�,Q��罜"%ʵ��)�Ǡ�Y%��h��N1����:BY$j_��m���OW����G�).�Ib��ܦ����2����q)W�����Z�]
�^�$�-���~Ir��vYި��+z��R�� �I�+����a:o<!��Hqo��Guo��ݺ���J� mP�gj�G֟Ȫ�7r{��b�fƿ
�J��x��{NWb���h~Â#������F�f���S�Qؒ���v����3({�^0�i�*��
�I��ڽ�sbEv��;�v��<�VYl-�X��)y��c/��^5~���������\g3�*��MQ��ݨ2����{	L��jr{����R�������=.|��3r �h]��XlxVHYEB    4089     e40�� �F�y� g3��K��@wzq0��#H�u����],�V`j���#4uv_��
s���ڋ��75K��H��fŲ�)i:�Xc[��=���{#7ETT�6I��꧕���դ����Pky�I�a��3ͯ����X7�ik�c�0L���5��>vt9� 3�����oD|�(���*�%\�#���Эp5"3�'h�Q��B����B4���C=޵DLp��kL5��GbE��JJ�8XE��aއ��^dss_�N*�-:Jʱ�5"��J	Tg[>�\a��낿� l"'%8g?+�@T;�0,�ӻ��JU{����!�C����	�
�d�5s��D��B�W]'|�A��Φ��� �H���6@3|�2dn�Gt!�?ynG�W�
�]���'�̼/oƶl��H]�CD� $tf<�bO�V�F뱸�ͫT|1�D�����i3��˜NH_���<��z�ň���+�H�Tx'c�H	���o�=�c�N���.��X��Ғ@Q+��������X��vX�:S5�Ĺ1�МsD/�jZ��p(U|<N�-�v��m[�qm���9y�	S�g.���U�3���
�٭��ʝ�Z"@�e�@��Gq vy��2n���@.�YvzC)����JC�[z���$�տz�?����5�H'���0yF,�:�#���~�<�>@���H���5�]�&����V�鍬w��3wl� ��ރX!o�P�״FjP� $�m���>�M©WZ���
��
#�y�ː����s�]fTX/�8֪�� !���������@e�EE~�uu/���/9�C{�42��AW��-(e
>�޽���<��s�ק��_٧�"2	I��lx��fm�@巊�� �1@� ���3fuC:���$�������Y{@`N���]U}>l7\���x���EKHL��N|�G��:S�1���Q����x)
Cޛ���гQ��)�z����?N�Ekm����=�m���E�ލ��?�/Xwr�~,s�O9�k�&�q�"8ro�� �j͎�u	1�������E�SU���ۆJ���T'7��m��1�Wx�h��-FNь
b����	�h�-��D\��a�����(M�g/)uͲ>u�W�3����á����T��ߗ�j ���Eiա>Ё'����mM�%|"�����.t���K��Z~�h�����`���2�ϗ��\���&v��c��/̷�1@�R6!��ዸ\�rͨTV�LN.cC��؉^�xH����!
�t�y�.I��g8i�"�܋F[�5�\�j�7�X��E�WS/�SZ�,���c2��6�����b���#���n}<kN���0h��ך*�	͙��o\�yOO�D0��0r|q�_a}"��Ϡ>�>R��S\|o���"��>ی�B�h<^'�KS���2��4<pPML8X�w��ȿ�f<��v ������U�~���.��:��dKy���7Pd���X1�a��nI��(߆�݋�o�1 �*V:�s�y��
l��dڏ���j32�t���8U��RI�n�wx��XQ�h�f��8�шK�z��{eH;��V=.;Ca���	��"���%RZ@qEvp���
�xD��o�x4��AT>�c��Z_J�~gH�޾-A��37�\��Qn�F�鏅��c5aw�e�~]u�Ɋl�C���4��[�Mg��Q��i��C��� /ؚ��~���(\�.���zd�#�m�a�ڪf��L���0����?r����q�-Ӹ��pW/�?E�.�R�V�~��|󓝠��LA��j.l�9�hOՙk`1��~��^MN%t�����g��-C̷S�ҙM�Nș9 H�%�D+ܱ N)+yU"Bcf�s�H�#����Q~M�e(�i<��hֆ��r4f>�}����p��y`n��,��S	���$G�1�6��'�jC��t��z����NJ��
��u���*���ib𷋉��\���͂�ájUU�"���Jg�0q.r�ݱy�
5�Q�@&�(u��׎;�TOGa0P5�km���HRu\�,��ۋe:�E'���v���D�A+Y�z@?K]]�a J���M�`���鞶>N̡'��N`xDf3}\!\�23���t��\|���g��lK]�?}���9��A���8�@��J�ShX�x6Uib{��p����W���9χ��q�e�d.	���v�$ ���3�B�i�3{��м@�\P
���7��_��8�C�A��a�t�U5�1!N2�@�:WW5Qg���l9�U���H]� ��m�	�Q�r3�N�nl����/j����m�v	�X���>|�{k�͔�x��yn����0��D|��Gx��d������?����MϽr��|�w�0��s���D씫>0���������)����Gf��O�hc�F��K����������jd����W(��9��y=���u����!�c֩9��������Tų�E)�կ���hLj�=�dȪϑ�xCix�*P���o���g��*�5 �S!�
�>�b�^	e�c8�~�?��r"P�����YWU�pN����*۱�s�\#�����Y��V��u
�C�O5���`h1������'�:�a��/-�]���x�!0\+,e����R'j�K�X>E�΄��5y�ȁ^�P# o�5���SԀ���v�%cyW�
N�7��Hﲃם�sVh�� Ճ�zm:�*��}׮�L]a��PWN;��v����FA:�%��j�n9$���^�Q���2����~O�VZ�%̛�*�?��-����5j,��֗L��jz����zJ*>g�9��m6�u^
�f���{�.��B�a.ۅ@t��Jƾt�&u�G[�:���}��V�D�5	b�|9X�-��n�Sv|��ٙL:�N2�)��>L|�v���p��3)�t����$�'���+�u�췄���=�9�zt6Zn�� �f��3?7,�	�n���A�T��b[��9|DQ�nE�ޛn�(]�e裬바��SLz51�EBM��ލ�fӖ�QEiߝ�o�:�;��G�ݦޝ�;�����9ٮϗ�i��8��om�hbg�vӨ�F�`H7�y�b�2��;�����;��"���/�0C��-WB��Jq�)o��kɎF��b��r)!�?DS��񭡘�����y0ԆȌ���'A�"��ߌ�������Y�jU�@�����q�
�7�I/" |��r�E���֑�>���|%��q�S!6�{��B�p���+�"�Z`j�����:0�C���hG��-xL�. �j�!�iH�5��?��Z�±�+ܭ�h$�Φ�2�7����f�l�]n�Ru�Sy��qu�p?D�- @��l�u�HԴ]2��H"�Ç��\�zl�5��iђ�q��̫	T��0��}����I!�r�B�O�B�z�S��֋��rC�Վ�Q�� xsd4y�x�}��L!-׮�_+�ۨėz�ʢ}��&��zX��|���[�{�(���yy9�El�i����.�:X