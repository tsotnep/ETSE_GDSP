XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������9G����:�q�̓h�vp���鑭����|��
�M��;��H0Q��$U����M=%����Goa�RW���'��"&���(�=|]1�~�[/���<e]�����Ҡ�{�������%�fj�篘�J�:��G/���Yh��R�*�~j�\8^dN��_�e�X��>`Ei
R����ZȮ��@��$���(o!V5,6�����|u��B��A��t`������9��q���l#�@�0aN�-�9�l��-oYmL箾��$辋K�J�W.��P��	Ų`���l��_ �NU��Ag�QC0Ύ��V�y
�&e�����{�f�-�gU,��·�x�X\�7�#d�Kx�Ţ�W������d�9򳜗C
$j���6�.+@��pH��f��-�;�˻���7��T���3 Ǝ.�;��yZ()��,N��&��}c;�^����*����yu��5-g��NO%)\��~��&�^���Lؔ�G}��~��D��B�II)w��[ć���B ]0)R�a�g��g{'�����O���SH_0�IԿ�_�)̆B�t���?^�`�qa���<~b�Qy�CGX���/K*?x��W#&��`�k�Ʉ$t��LQ̌b���'y2��A;�r�����Y��>ĉ}��|b����i	�y v�(l��a���%������f��j���V�\�n��T�A��b�e������>�aŊ���[�YP�,�XlxVHYEB    fa00    2470��kGp�*s;]��ċ�*�!�Uw}�=�����.��=���m�7�g2 �ָ���W�
��ڹ�
�}��)��ޫ�1�zyظ���il����!�1h�s�8>%����[x.Ix}N�n*��j������R��<��ލ�
�ٮ�>U�ʇ��e�t����Et<=�m�*@�������S=(o>��g��T��	�r*�x����v����;9V�y�"�x�9�A4#_�
���X���Q��)
�<�+�@fӠE��vp�r[Ѳ?��V�)-Ƹ��vX��	��!�n�:#l8b�_�6�Ac���Vs���!h��#�!+#�E��ǘ�x�gq�͐x��X��j,�ʻ����T�pB�n|�n�H��U�5�L8hP6P�^�w'Z��F��Zc�-ǁ�	iC���vQ����<�r�ޅ���t%��mQY�M"L$���1x��5p��#�e��7j�.�b���i���� ���抉F�*�����[�+�4`���N��V�phoKTV�%w!�b��]����i(�+r� ;G�'�-	���)c,�g�Q�8~�V��_t�C���K��,���x��L>Ƀ��وez���%��7�rG
�}��uϢ���o�{���+�XY���`b%UC�'d���p��e%Z��]���Q���N���Q�=a�p�>p�_��%������v�t��"	�/������S߿��6��o<��-9�'Ğ��.����Ai��0�/\����7�eؔ֍�C�g&��s�9��K	t88�R}?s*ļ"`��-��wܜ�5d-z�)�U��6���?ybbX�k�<����F�c'o�������v�����d�`x�뤔,�!6�f���b�TYGtR�E��^�K6-G�NT��a����EhշN+��Ub�L{���F���G_ucJq�t���;��e	@�D,�kN�ܗI��TĢ0篃��"�����M^|\���5���<�bP˹��fBƔ-���6g����E����9&�"C��%k�C#�d�eΏ�I�j�V�'��AU�}
�S�[��I2��T�fN�v��G�u�7�>�}A>F�D_Rj�
^��Q~��
OSX�k��{ ~��~�ɬ��`~KI	$:Nu#��s����Q*�2����e���b�N�D��(�74'�%B�d7���K)r�	ܽ��q��}����bc�,��0;��^c�����b��¦0w�KӡD�Ϥ{OT�Bh�֨&�0u��U�^���p`�%}�F��1|��lff���i�:8��f��-�կ/���X�ĩ�iM��?�)�E-�Eq�n�Н�3�;�X��z.���E�`vj}��>�[�J����v $�2��Ys\�f�c��К�$G��Û�{2(&0�g��[a��C#�v�쵆YJ(�$���K@n�@Ca��|�O�>��\e"m�Ύ�L#�c\���,�������h_�$�栞H�����b�v�i�~�9f`Z
A`ƥXVTJ�V�ٜ'lhC�!��/<@*Ӧ�q�E�2R��v�O#M����m[⳻�%^h|����[b- \7S�>���U�)�W��!nMW�E���������Y8*"n��<��t�)����F���3�mW��� �~%��)����y԰ep`E��KPk�ɥ�JBH���g���%��-�Xg��� �������N�JK(���߀��[�eZ�˛+�ÿ�ah���UjZ�K�(�p���iKBj�PO�
�\��Z�v��I]��k]�,�q|���Dz@��׸�zɐ�B=�4�Ѽ����$���^��"u�`�vǚ2fX�$y�F�7��	��ߡMs���I)�������CQS�����U�O�k-��Q3*L��&B/����(�n�R�IOk��{CH��vr����u2����h��#�������|@&��|����3�����qY
�{���Ƌ���^�N�9.��R9���O���<L�p�o�F�ѱ��ߪ�a�J'��c�
Ҹ���9����/�� �fd�Ɏ�V�E�Ģޅ��T���l��'u�
�B?c8��a�A@'ns�7�J;�b8�=�R�ZuǇ�"�ڧ�,�$ȡi�� ⿰�����!�������Jv4 �ql��6W3���B\"�+ec�N��8�z���$N����D��B�?M����bp
�u	���ŧ}R�Ƣ]�є`�hͩ(�զ�7�:�O*׫���:J�!̑k.�$�y`lB�(5w����HM��>�ώ�a4TAnj�[k�Yu��b��bf]/X�6/�xg�E��ՃZ1C�*�D]�_}aUw���P�z�&� �5+��'��ż�Hݕ�x�#�xT���@�{e�jPQ��Q#�8�q�loh�.W��
*�	�h���>ejM	��A� ��� A�F~�A9nQi�{Y|7QKJE�XI�"+y�(�Lk��f[�=�4<+|���3�B ��\���>K��^���ϧ*���w}�<��yvQ��\��Jk���X$n� d�G��KD�$B���%��w��u>�*��'z�����61�n�t�<9C{�|�w��$��r�^�a��L��.�O��S�3��g>s�F��%8���?:4ߊ|�P�r7�h����B7�=��8_x��L�`f�Wg҆���A��8���k#Ї���7��׻pzsA��_OH����+[[eВ�#�j'���������q�h��,.��ڋ�u`��b2��\?�Q�Q��b��oG�T��V_a�|�h,/���7�Bk;��R��T �CvCu�V}欮Б�+��'��E�['MUl��o�GA�9N��O��s^�����{�,kS�a�ʞ~[�z�]
1W�;��Nl��V�s�&��ޜcw�ـ���$i}�Kf<x��K2�.��UV���G8wڱZ_u�ʯ���z�h��VL��,��Z���9�n�ތ�nOш�.�3�8�4�� :T������r+'�oJ��¤���^���/�ǥ����w�7:BhK��{H�ؽ��ȟ��	������/�N~��^d!�u�E?Luж�������WJ�n�~��syF�������?���h�7��I��j�o)[�:#ɭ�����O@Y�"ˍ9D�n~�4	�
tɊN�������Dj��kl�|��G����i�p�^�m�F!h���q�w&�]1�Ԡ��@	b+*�z���_�I��e���Lk��_ei��d�^�t�����u�0�-�\�2�R��w��q�L����ڭP}7�u{"�q�#�
��?�@nH��x�$я�U�Ov��r��<��I��&��!�p_�/݈�=49x7�9}w�`�L#,�<!lѾ������L�5���]����-N�pK��+��ra������&u~u�2�?�?������b�i��ܱ�S���,j��j�W�9o���n�s4�h6�6[yӑ�>����|Q^�nG(C������i���|����� Z�L|�G��e�B�mNyV���aƖ3d���8�s���t5uLr�g�AoK�~��k��̿q�[�	A�su�qO6��d�)&T�bI�G��cx'�?���V��ącƻ�H�b+a&Ϊ�˖d2Rt��RQ��D��;N������
�q̜��b>�)_ky̥p7�(6ձ�2���Y��� ��q'W��B�`#@Q���{�.-�0ӂ/5��u�%m����`*T�;�lc�0H��_t���߬(�\���OȲ\>@
�oﻻ�l�=¶5@ҧ��H�G*���q�%p$>��4���ƶ1�z$r�_K����:f�H?ʈ�P�)@t��P�G���Ɵ<�7�c��$���1p�$v�����ھ��~foE'P�G]cCx:sih�C~��]d+�y�=�xN@z.�F&��c���1��6YIx����C3�`Pp��(Q�]�Cn',�/7Z�{?C��3+t��k�)��'ft6�O��oD�7_5�p"�|��Ȕ�� ����]6{�N	:�Wv̂sk��O�#/�	���2�y��6�a[�Ћ��t>�M��{#��9��P�nWi'��򻄧ӿB&���Q��|Z�9^Gn�ۤ���]�qf=�qM�d����
tMJ6/b�e"��N e����s>�wE����kl��[��&��_�â��@ǡ��Z��̓Xe<�œ�0M�8�!&.!�6�*߆����[�xx��M�xG��/w�}ʑp�Ɩ�c�u�tX��z�����8t�4n��wi"�&6#߻Z��T�d��!��N+0\��H�6o���E6�)�9<'
��M3tǮ�Yq����z+�����α�kB d;�6���[�d��6�AE�U�"Ş�M�g̴7�b�i�/]Ʀޫ�Ed���@H]Ɵ��?�%ec���!��O簸v��.�s���/����w ��h�2ʱ�x:�Y-�k{�T�BA���KqY��.yez�n:�&�w�Q�YcZoJ)��Rj���J�2�(.�e&���4Uwq�:� ��pk����!�1N�2���;�n�b�pPO���D���)u� ~�
U�ؑ }�)lqf��T�׀���Io
���a�F[�!S��$�a}���؏�Hp�`����i���?�yv�L1���I� ,��L������!�j��L#w�hF��3e�r�I�!j.&�ٮd
����#�B=&�s�FN���{��dy�)��̵9[%�T-�:h�Ym�`QO��R��W��yg ��p��ҳ�u�,4���\5��o{ׄ�Y����>\e|����(��;!�*����I]]����*�t�֔�� �u·u��σq;�蒺T�PAr�B_��д>��$����[�$i�(L�/�/��;|�<FE4�
�=%=�s������f�w�
�����A����1y�
��
�n�E�ݟIT���Σ"����譤+��'��� iQ�"0��h(:��Z�ö����:qxj�ta%�{�N!;���%��8�w�) }�
�9�0�o���C�N5F�΋�#o��K#B��A�Kc',Pe��q�@�����>����҃��6�����xj&&��ʺ��,-)���g��g:4�~�]�ϭ@��Ǖ�r;�����a�n�L�'�lul�c�d�7i?�i�7�!���\J�W�5�A�Gq7���pOY��9�z�y2�y���C㌾	�8��F�0^G����cd�,��:,F>��r~��iYr
�jx���
��2yV�%bpI�	�e[֡�0�j��)���3Z9e�wv#\����i�����t�Cs�'`3����4�n?pg��@���y ���W����sr�X=jm���kOJ�ϭ��_d��P�b��܎sӹ)B�5f���`H�Hl��F��I����𵨤�&�����]ƙ�#A���ϰ2��02Ӷ���8�����OzYm�|f�������2�nh�ג��X����D��?A1����LF�1�)����JI�����N���E3�0�,�y��^�_F�X��j�B�O\��3/�ã�ZJ?�]
vP1]Rn�^��A��.Qi	�d�N,�m���e��1����4B����sy$��;�c"a]@�O���dθh��eC��\��Q�a�$��IO@���;T��}ף��H��2��g�y����R.����=��o*��У^�'��U�ۺ��#�ۣ���z��<��q�{$���������aJb�U���CG;ase�p�S׮��$��+'7^��f����)����K�zR ��:��X�[J�s�dL�Q�ɷ�C[�ս��Ȩ�L����<��Xd�2��Ѥ1;�Y�����-���o}9�Sүy��������T�Y��+�k:X�z�\s5ƛ��¨��/�&�,)Ek����%1砒�/�x��P���$I��2���S�e����.�z�gVY��a-"a5ʇG֩�@P3��P�5ڪ���31��o�y�iw?"d�q�!�/1��B�ջ�e���،z�}懶Z^�����`{����o'W�o*��ˁ��L��ўwxݼv���؁5^���lo�O����/��:���Eͪ�+4��-uF���g���1{=�R��b�i���ܫ�㐅��_�p4��GG�-T0�V��~��S��p�����^&��##���j�IV���l�����C�c�P�!��o������%/�,�Y?�w'�2۰4g6@��*q�܆������yţ������Ў�(4��Ͱ�J��q��J5�%Hdஅg�:i�ip1"�+����(��,{�77��{�dKU��燎�o�%6v��Bmn�5S�~����紟��Sy��D�����@XY(�Wo�C>8ī��@:��`��
����*{��M���]��y�"�_�φV������zkjL4NާRT&���Ht�I-\��&H���M��O�,T�>H������5X��8�誾�G�qQ�x�IcUë�"� {�� �C�~�sI9M��vZ��X�<�L~�:;::���ЃD�%������.���h�><[��ETT�ċ4ٶ������烍���JU��x|O��(
`��ZX�A��X�Θ
V�9���Q_�����]m����)%�=�������ƅL������~���Y�����z �$`��f���q^]խL�.��tI��0�Q�T0�4`��txr�-i��
���h3�E���s?٩��w�M�l�41�Fw��YK�s���3i<Q�]�:_����f	k:G{F�D��"f�̊�Y#���ʯ��E[�Zv;]�=T4�tR$�ݺZ)�2fdn��'J�	�@b����u�T!��6��un�SLc�ʞB�����y��N+�~5��u���iݣ+�$��m$�;I=פ���Xɩ�fJ}^��k�����,ך��;���R�Es�O_&=���
"79���g��t�N�NJ$������<�fPR�Ǡ��u�T�6����=��0HB��D�ʊ/M���X��xo��?B������l�+�z��
4¨h5�J���B��n]\9�-�!<I�Z��&�V��h���e�h��X;����1��a�?/�s���F3�~Ns�F��з��[�g���ʤ(�����vE���X'�h��wbFp�j�aV�K^{��rd�|��'a�>P��x��y��=� ���5z���LZ&o�T��N(�#��P�ar�*��|�3�rP2��b5AH�҇:�4�;��o���+RO-��(m~"�u�� ��$>!�d�>����d�MK4�"d�}d��Jy��_í�>{�L4\�4��8꼐�U�
w�T��R�:��)�I颰������q=�hŪ�:�ݝ�Ah_Xr�[şj��8�S���d��w~WWL1)da�OH�~�=&d��9�!o�w����yy֢�d=y���=A�V�w���i�!���VY���*y���k[������[����v��/(Z^�����BK����X�+"�w���.k�G̠M �������B�߅�����#]Iq��ZR��;���3^��� i*�V#�U�6S���;t�?vp�E$^ř�ac/��p���p��X��l���fD��s����~��5ŀ"˟��K-��7����%w�/�0�>��a����f]}O�?S�Mj���o���RR��
^`��"|$���$�r2�8�c�W���o��'#+�Γ�RP��ܯ3۔.qͫ�"�r�:�'F�pn�����n�����U��_%�ᄁ��'�Y��<c�|,��gjq;Z�s9�3��A!lj���n������uwƘ6�h��^Q:M���S>��TK:����b�0���&U�zx����] R4�rp��aD�*��.D���4y�rj��&.��4�2�_螚`�g��cQ�njh�s�����@5ò��-
VW�'�h+�KȖqH��8.���S�5���EZ�<�v�f���Mq(=e�O��~��\!���Qc|����&�LN�f�1�Tl�2h�vV�����O��?Vc\��u*(;�~>DK���l*qn�K�&�"�Sn�|:��.���o5�f��N�#�MCTѡ��p~c�sm�m�����z%j�\�5M��h�O�ad�y.�Rj	��m�ЗՁ�!'�|�V8& ��y���(�x�t��ߺhsq�9�L��������xX��{�YM�|�ѝG�dn��&����ȳX�4�i�m�"A�FUn((&$�?� 1����	���8y�����y��ſDU�,�,��9)9�5$a�[��P��Q��EF�(One8mv)�^�1kn]�k	(�JS��gV����ٕ�6�:7k`�C�g�Xfb`\GؿK��{������NA���^Y�W��PuwezܤR[5��R�$~�9Ԟh�4u�m��Tm�cD�&�d@ʀA3zsJ���#�o��p���	��q�`�﴾	��q^��$��V���-��v���(w�@���"y��[}���4��k�O"�<f��_P�/�Gsayq$�v�������N�v��(�}Pn9ZT����s�ɿ�c��t��Y@�����jo�"�[�xr�[N�����̛��� �J/���?Q#DU�h������X��kp$xl�X�h��_Ì$m��B��&b�����$ۀ
����B��L1����3
�T3��`�:�N�m��9*?+8~W�{qMF�lPŕOѥD�(`_	�6�>6� �$视NqR�1��_�E���!A�C9�֨���1f^1�+�t�S봣�-t!6���a�c���o�P�'��[��!ܕ�K�[�[�/�
��\��9���CXa'�8������L[txX�<��2�j<qp1z��Yq�$~b��\�UWA]�����a#�5g�)�ˎE`��e�tXݪ�v�piP�H�~Ro�n���'��f}M��P ���1����.^�s<DBA���Z؂A� c�ԏ��GLH:�Š�҉�-�r�>�8��o�e�Ŏ�4}Ն��(��봩��<pޚQ�,��q�j�(�����1��O�8�aw�&��~�̀��h36杉(�w�n�Z
���'*��U~��J�d,����Q�����S<ԧ��ָ���]�����l��4�  �JX�@oXlxVHYEB    fa00    1b30m������]B��qw�Z���
�͟�#�[@P*6��Qe���`��!D���?�Q������nkK�� P�;�����
^d��BTc#h��S���F�͠�
�̕�mݯg.�f��D_z�X��
+�G��%�s�����p�pS;!"GO�gS����u�����.���%F�w�K�����f�7'LP7]i��W67�4��d(R���m2Ĩ!��oi" m�����2�0j���, X6�c;���� ACY'8�]ُ�c��`H��)�{�5ke��b1��);(!��9�+���~ZvO:�zv\ɦ#r�F<�4�}h˵�̐3�p锃�-���A�P��?�����m-T�VF�qu�ɚC�Ac��Oʭrx�l�ޢ��ߠ�@L@��?#T_/o;�*G��ݰH"�6�"�,���� �
�s
�}D�y�R�ڹ�7����qk���a��t�?ʥ����!F]�$�)���S�
K�}㍾l����s��j��-�}!dIl0�f��J.���lIoL���s��m�SN +ziҏ�X�6")0�� )�nvRA����|�v�?�q>���KÕ�R>i9Xa?ӟ�m��;˚2,��+���顃�z؏ =��uxǗ[/�,:h�ޅ
f���],���~0�v�OA?�k�l�6s�*XȐC�M|�M.hӑ���w��.I ���ZB`jSdqW^�<�Y�.p�W8��\�F�����=tA?AuvnS�_u[����c�����ƅj?C=}M���3S���5�XM�WG?i
.��
��e�d��̆_�Pھ������#8�e�^���w7w���2�+� �6H��]̀�*�l�T��q���݈Y�.`��'�6����x~��5�?��͑<�G�ޗ�$*�E�mq{�-�BkxuJ�?q��[�y��yq��.�8�xnh[X-g�E���O�[�6�칺���x%�V�k���!ݻ%��^��*�������[/'��5�@�{?�����N�_P�h�gl�L��wԮ�]@���j��nВ�ı�ş��D���+����@��@�/��:�kUu1#�*�}��d�}�/Dt=�!6R��Ls�v(�� Og�h���e[wW)n%�A&r?�>��
=��$������3��9�ߍ�<���P乍@�#˥����fXl��khPc40㏣'r��D�Ⱦp�7H��*UY�[����H����nsx.̴�]^_u�n?=�<���^*��??���'��kz�D��K�g����z�<E�F8�_���ڂ��D4$&�Xl��z)�w����m�����'J�$��-�֢�F%��;���-7�.3�$hdD�Ŗ-�f$��00gvc��p@�,�+�l <^��v���ȩ�6-�j|J����t)�W5gr=��Θi+ھ�?��.Vl���)ϒ�M���R��YM��p����x.7=�P�������de	��X"R�<��@n�Tʄ�n>2���ڪ#z��Q2�������).ñLjI_��3b+yJ��<�ҍ��(��Y�ұ2n�Nm�q�l�H��no�ϲҧ�o(|�.����[T_%#�!��	.�٠����������A��]���z��%�樦<s"�N\[��Y9��=!��`0+����{ݿ���cڡ�\[�u�"D��1�������f5r�K�v�j��t��������sD� ���3�b5��0ׁ�)��~(L�K���.��5\6&���,�x;fEht����Y����	������S��+e������ӟHƑ�x���w]B���kF�IX�Su��!:�[
=Ro�M��|�⦸�ٙte5�:�^g�b�����-;59#�㡼��c�4dh��D#f�Y��:=J���i�U�fY� J.G������"��*����;���dM�v��tu~Q::OD���v��d1�h�a�B�T��?��ު �	�J��M��u��%�}2ɽ�g�"��n_3�T5�^��IV3����6J�Խ�&��'\�X��,F5��v��S�K�>8�zT{j���(nԛ�v;$�g2a�2�U;Rs�ݛ��'C+c߱B/w<�VV�����خle7�Y'����˿�����;��Ha��$��8U�?AkH-%e*�^|�����q)�\N����|��w�)���v|�HsK��}��|)��K�����IF���(�E&�G'��#�Z�1�v҇�Y=B=pU]��!�T%&_\Օ�V4�괫L���*�)fA��}����w542�]ᗳ��F�EĴhH6+��C�@ru�v�F��&��N�x�0z��L�RiF�)LW�U�>9&g[�ʔ��=���ߋݣfu�Z�V�,~���L%Ϋޟ�7v6�'���G��Mu��j,��I�� �5/����O��sD�=��-���U��YV��T��6�������bFa�&:�M�;7�S59%���Q���r ˪�x��hu�Em�@�(�bk4���g�.������J+�쇑38�/֣�D���� �+�}9���Do�����&��Q�f�
�b.3Q}�n��d�?D�\�T/��YO9�W۷ ~�LS��s����{Z\��$$ˀ�|5p}��!e�Ό���j���w:{}�{]\[��gmR�0T"�Vi���;��bm�?5t^T ���:S�s��PB�*D*䌹��u$סoU�>������$����H��9#��ؤ�3X_̒������O2��Z���k��~9N+d��z��+#�i�� k���;$Z�~�;��P�"�{�
��^g��1�w��c7x\[y�K��=�F?S�p�PS#���_�t�/Wa�v��Lr�Ugp����U	![\��U����V���������kc��QM`�]tL������Ã�n�!����d�2�je���V�=^�NW��X�?Q<0.���'�H�\�]���!�� ��Y�&7�����F�W(�2s*N�Ӷg�[i�ܣ�,25i�zZd�@��zц���H�6�����HDQ�v�}�ھ�YOP��h"��f���=:��� B���&?,�*�J�OF����r�ɇ���U��@k\]�i�Sq<	�%����L �`�(l	�2N�;=��{����*:����!��9�/1� ��-�[IH����:�P+�$\Gg�&颞���Z7 ����oAMђئ�te׮�#�סZK�{Us�5�3*�g�@1g:FB0�)�'y<J� ��� �������<�b��o����B?�q�i��o:���Z6��^&1��#~
J�w47�w�;�$F����7���Z�w���L�0�Pki�K?��D��'�Kk>蝕�XA��_���Gt=}?N�%;޴P�Ml|\X���\�ϗ���'��O�����p�dف�+	�"(N�	G�j�e�#�ZL��7A�m����s��j�9E�ӉO��wӾ�eBW���	���s�9����� ><�c";j2	3n��<B�ԍ_�]�^U/��-��t6{s���\-�C�sĸW^�:��V�A/�@�c�;H���^O���<2��-��ɁuU�f�e�|�wKV��S���U |N#��-��;F32V��Y(��L/���$��#�yZa,vWvd����P�Q�&�PV��Q	Z�{����#sB/3Y����rgBz���NL���/�X�W'�GQ
f�]�g��a�]�]W����-�B��(	[s�g���qK�\͞@�%�*������eYl�x�Y>b]���f	��%�[b�-nܒ���`�Y�#��Ԕ��L��G�Hp�@V.�����۫yY|d����UJy�%��/y����%C��e�r�Pcv�~�U�yw��lkЀ�J��;�6"��M�=�4�1�8�7��7i3ͷSI����)����S�P��Z�a�
u�q�����ڣh�G$��;��M
��dR�˪G�Ow��Z�`��MQ0�R]+��eFͲܹ�q	�cUN*˦�~]���~�rX���;3|������2ko�,�
��b������'� �8����_��{���b��֖!�PMf�Ł\�l"�S�ف�l����yȕS�բ\����?���J��^�D*��K���%ĶV*���Z;1�,:�����Z>$�PXt���!�D��Ի�lٴe({��d-M0O�c�}�Tf�������w�>#��ڛ�K���i��5�Ę���(TҬ�8ڑLw(�L�{?���]�Kh�'����̈́����Rq�1AҰYoZʜ�_��=Ӗ�H��o�}S<����e :�	�5���*�!÷#�8���_���k���}�w�-~0���^�)�krcl���]s�L��iQ[����KaD��I����5�f��cf!��������-�L����!��=ӟ	y9	���}ۃ9E��;��PԦFa�
٤G0A�^crK��f?�Eb����d�:5�o��?�^�t��ۆ^�������o�]<5�S 	*bǌ=��3��髎� vV����"���t��_�b�Mq�g��4sQe�1ܡ���5%~�~�/��Z�jE�5�/0�^���0��lL��RNWoB��NV8�P5%�AQ����%ǲ	% Y�l5�VY��\�.�PA;����6.�͟X��Z 3�X���Zc�؍�L��J���0��:�qG�����}���¬�j�
Y�B	.�<4�`R�!���-h�BB�{��}�q'�f��wF95��q4�������D��`&�y5s�.lӛ g-��(a���[��'a�ٽ5.����'?V��=?e�#ɪ +��UH�	̉���=��5*��7�-�������e�~�^N�R�D�B�o�|5�~1�Jlxcs ��PJ4�������P0������\�\��]� ��W}V��b�>WQ�����
���Uc�^��%�'�+g��v���k�tv>�D�x���נ"6�gHo-,��g��Y�,�j�quD��Fl�~]��6Z���5x�!}��W���d��wWb���g���$y�U"O�jk4q�)���9j¢.��25̯(��I�<7e�v|؍��/����#������GT�*a�(�l��l(�K�Qla���HXW[���G�J�#�g�ިbj���X1 �p��@�D#�JC��nHc��1��͢:�^���(o��t
�f��d�����H H���haA�t�u�W�w�0�E�"�:�zvE���C1Vabu1!11.. ��ǟ�"� J�ӱ�ME��P��bU��!#���2�?܌mF�A��� _7�<��P�&N\U#T2��!�/c|�Yc�A�2D��Lw�&�F�b@!�%@'";MXD��)��E)�3t�J��oQ�)�ѤxH���8�T�^�(W��U!.u�uV�4���`��Y��:�t��ޒy��Fh�߶-3������2AgX���-�}�ֻwz�-)���IH{���p�Z��;Y<��5'k �sr�bYd�7�� XVEk%�o4����@��3��n?��#��i�����/i`��9
ϖ9�"��*�Ur�+��ʾ��cMfj��z��k���_j�Fj!:��?�Ɛp�3������iylu'�������=곽�KOEM�a�gB���$�#q��h�&���&U�Y����3�L��W6חm�4��LJ��P3�#�Mm38%#T`���R}��,�������%����ܾ�| ���,?�ޑ�R�̓ua��Ao��U�G�F���+J��KLp*=���,�!��τIsXv�����31U/��| ߆���9�ôVZ9Ey���$b�H��a�_��#����	��9�#zui��C\9T���g��`>	�GO�Mu�6�-ǉ9�U�ͥ��*&"�f;k�C�kj��\u<��}�� �Hny��*��&�RԠ=��X�Ǉ2U�˲^.�H��<'&P���-Nr�5�&�0�
��g�A��I���k�,T0���(��wG��
Q��$����!�>�ǧY9�|��A�~��Uo�D��l��	 ל�^FR0� ��ZI}z-�\߆���}RM�NS��7��ws������(��8�~��\9�=��%�Z�ˡ�d}��)�\�QNE:�/�+jM���H�U�u���M'�g��{��~�g��"0U��퓛�uj��8����-�� n&ȲYoA�A�x���@3��խo7_��"�-��<:��D�T}�9�����mN�m�Ef�R��z7���(W�nwJ�dF�#8�i}���A@IN2/�F�T�L`:���pwo��sҽ�y�1��?�ြ�ۣ{�B�b �J���)���r_��1=ã�����2Ϛ�4,��B�v��]�: o�,UA�&����	]��f#�0kT�'��u�GJe���ݹЍ��_�5V�X❃��xr>s&���SpJrRn9U�a��R��Y�$�`�h`|'�$O���6�3�j5
����*���]qp���Xql�.�
������:�{�9;y3a�+��W���=ט�aof��+�:�tjCaE�]y�q�
�DNN���^.pd���)��9�Ƒ��l�&^_�C��'78���Oy�O�v��L��w��f�����&h�L/"_��ݓ�|q���W��]��R~`C{)�HIy�Fw�K\��{���{t���L�
w�Y�R�W��b@kU��;z�B�U�=.~�\�%��E����'����,�DI�j)�@��>-��:�^8�@���7p�4���@��XlxVHYEB    fa00    1950�A��,5�eெ��+=�-NuE�ӳ��"װg��a��x�6k������Mn%��v��D	���W��p�T�6{cE���Qv�?�w�*c�+�'�(���m��Z�N�h�$���@Gk-�����0���m���S[V钛K�;����e�Ah]$P�h�򉱹�y�����M���b��e��A��҃6#����@�7��D4Ͷy�М}����`A����fCE^|8O���d��ߵ�}���r7���^��7�(�\�D���{整���߀�"1,z��I}M�]��x�N�<�6&�J;T�Y��'�Ac�0�H��f��uyk����xғխ�.��T$@eD�x�Ay@PG�y���u���L��~(r����wDonb�-�2��ͻ�G����w��Y�Gԕ �[Ft����?�}��~Xxy�	�)+tg�:���>��R��&q������t��n��
�\�eVI	��Yq��\,46SU֗3X2���l�p��5�epR�\<���BUDF~��y��!�ί��K�R�dTv=I(�sz�����Z7%��BJ*�Xd�����lW�3E����:�Îޘ�X�(5�BY/4ǋb�����6�rx�4`���J=Q���}Z.��;�µ]N ����H�mqs�@���z7�u�O0���LTS�ք�/�l�u��YKC�9�e�,�D�#�z�+��'�cΊ���x����2�f�w���U��s~^�{�r^�骐)���x��c�Q��W������r_��Όiق�ӗ�=mg±Qm��_�;d�Q����WR90	��" ��>��2g��;�j�Eɕ�c��r�m-�j�"��dl�A0ݦ5)
�ˋE��2�Lp+d*]L���'��БX�?��|�A�w�ʟ�Y�mum�N���aX���4�z�΁�S� �N�I䰌�"�@�*��P�&v}�,�����y�נ��"W}E*R�9�-�A��U��V��4�XR��^@�iE0Y �+�\��t�Z�7s�\�%�����S�~7��Z��gM*KW:�l٨���.��^��v.`^�sqH�ʥ/m��j�[v�
j�O��b�B�s|��:���f��r�_�EmHN�}1�0�p��c�X_�p8�� �Wz��X�5�4�����'y+�\If�j����Sbt���8̯pH��������X��0��V�?G�zac��b;��?]�z>ܷt�����ĸ��,|��B�=�d���D�Pf=� 
����^���=c���"��,�\KJsp�g{�J!���h��%���z��D�m���[�Q��sa��U�-/	|z:�R%HE��T�c�p}�L������.��t]0_��e�I.���ͦ}ܡ����~V��&^��RW.����
�w_�[�R�e������ȥ(:�y�l}S�f��>�K&��`{D�[�r��&��ݯ�"��~��g���B�7$��Dud��$�Op�
=�Zd{����
�㡒kE����<�utf�[�K0�4�X{���K�&�+�ܼ�7^��V�:�<���j�^��2B\�"twNl��!$�����V��H�V�h�z��_W�E��ḟ4�=��r9$e�� Xo�^\�v�9�(���u!��/��f�.Юf��6`'���?�{�M̀����<Bl�]�<y򶝁��g��LB�ׄz���@5ؑ3i=��Z҈\���깫�K(Q���G+�S)���a�E6�&u�K@�>'3[E��N�/m��X��t�BF('Z�
H���d7���t�����L7��jQЋ��t�内��$�Əكf)���cS����Y�b���*bֱW�V��}<͋ۄahAv�N$"�2p������n�Y�A��,&�h6t�)��O�'˶��%U��
�H�t)�]w���p��eMs����`4D�{x�_G����!n���4��*
��:4B�<���Pq-�����釻�nz�XU�����ʔ�͡���4X!eݢx�v���k�}"���)H:�� ɓ�@ky��e�{*����(+a�q�Ҡ��3��0:� �+�Wa�<%l|�F׸�;^���H/���LI�w��nҺ�e�i�t�X�\Ϟ�{|e�°d�T�Ýel�k���`���f�58E��XH�\�KqN����:�oI 
�j���ekQK�Vd&K96�r"��ͩ��"��e�,8��Q\�>��]�ay!�
U�O(�u8ψ�wĽ�RȖB�lL�J⤊����H/ȹ\�������г(�잵�7��V�G����M�cg���:FŒ�+)vU�F�Smh{�Q��$�W���ӌ���d���b�PQ�Nd8<�
P�TTT���0��LO\��J���r6�s2�
2�ت�~�
hA�mZ�d4�GF��@M=�y���LP��T ����Rχ�(�ЂxE��	�J!c�+r�����[��`�)����G�EO�3��ku%�J��J��l�RKL0��e3�lw��jN����uӃ��O��@�GZ��Ō d�������lo���p�����??ٶ��\&g�$1�~9�@�2��&&푳�T1*ה1 t��:��$p�U�.���	� 3���/7�~�p�i��ln��\9v}��d�10n��z��r�N��S�� �οƁ(C[�'�sɻ�O4���,,�.�*^^(�9lg�b�#Y���*h#�z{9�c�G������~�i�B p`�v�p4G5*��b*�wQp�N��7'�����bb�E�=�f�hrV�ɚ���(ˌ�,����8s�9��,����J�em�A�n�v���K�dC����R�x�I	x�*��h�A��]�p����6��͖��4�ho�V�9g�%#���(O!��r�Bn�6j��v:��3�ۦv��.���=�4̼�:���x�8C��ucΜ;�Л�DQ�J�F�Ix.��f�1"J�%;ܚE�V�=�̚����_�-9�S�H/h0{#uZ�a�d�^���d�o~���f�A*��3����v-�Jnο�/��+�RRH�<mGЬ�=Xm�)+oι�Vc7��-gW��A== �	���?_{�#5�h��#%��ע-�xƙ�q���w�y���[-L+�dP�!p{Y�D��u���Kx2��Oh�ф��%���?�p��'�!�Uu�!��Ws�a�(�Iq9�z�|����,]*��2��,L�*F�)�<�̨��ɢ>�@�w�f�������b_7��H�����AɨT��Tn��)w^�6�\�f S6`�Q"�c��HT��\�s(]��|���~D�@{���S��03�PA7�@�(�/#W�:�J)�إC�L=��"b�KUI�x���"�c��4[��U��[�S��'uC��ÀA@�0p�}ٌ��H^a̱lL^��౸���6����M��:���;���d�)М���P֕�o(��r�(m�kC�|e����S��0�&ÒT�%l�
��b�tg��5~�8���$oǀ*1j4#���3V��J6��v�,8F�)�坲G����Pe]�#�'�*d؏�#�c~�����b�{ �F�Wq�#�
b�ޓR�n��`(�����G���,a��;���:雔)�؝ʨ� B�,4D1�q�����ft��DRb[�u�p`<+�By�Y&p�.�&=<=� �R�78x�
U��.���S�*�f�$]�o��ij&��O��(t����u���;��;���T��n�y�+p�� Ô�����9�� Q �Z&��>�%�m����B=xa��9��ײM���[d�ǆ&��i�{Z�X�w���U)@�R��h=�����o�ܜ�B(����̏D����-94�����.x��,*d�Vs�'��W�(s�ڝ��C���*�#�v����'3�N�7��6q��$P6P��t���M�gN�#Y�7��C�MBv�O�\_|����kʃ���+��!/�n,Y8���[��Ӿ7Sl�φ����]'�o���{�e�}:S5�r�v��m[�������ޭ@��J�E����i����d\	�)���^���h>^���v����ň�Z���qӊ�T�{~ZpQ`��:[�hc�2c��'�ʢ���`fV�B��h��� ���/y��$���g��Q	~�@��NI�*TY[�K� ��Z,��J�}��cX�	X_N�S�a��7Tcli���0Ｅ��2FmP�� ��7��'�!�a�N�ω�m��b��{/���K�¦�R�+���ht�]�����M����cq�À�{B�z��eϱ�k,[x �@a��N��~���y�)X��&�N2i2=�0,J�{��mu���V�DwN8�>��9�ڬr�_BG�,��&��I|~�v��oE�����d:�J��I��ĺ�5O67��-]��X�:NO�#j�T2SL]31�w��1��9U� x�u�R�D�Cnwb0�p6�,и����Q�o�Pʻ��S�7��u\S���&iz�lz:��TQ���7�l�	;�T���gZ
%8ӷ3��~��H��D+�Q�� -X��ò�m�r��Of�����:����ٷ5X� k�CӾ��9=��w�/ò���?c<+���J�N��R#��Ts	���A��x�h�cEouZO�ŷ�I�A��b��}��vU���M�����^9��!aa܍�����j:�=,�"�c�`A�,����ʽGu�r�թ�%�[D/�m��H-j�x�1����_�t�+sւ�_j!�5��[�uH���gd�R����c��m�FK��9�ػ�{� �ZK���7 �(�TVr��9j5�\��	��2��R_҈�M-\�K�J���|�4�����ο^\M���i�]
��)��9�ݖI,�-�ϲ�#���W֟�jd�Gp	 ����)L�(4$�o��`��/��N����ߕy�y�@@q`3���v�U��Bz���L��%�9aq��rW�n�1��.3�Ǧ�W��^���?zҿ!#�o%��)�h��N���/����{���!PS�&������Z� 	I�t�T���g�A �%ǋ���v)�#%�����4,U���xޮ5�_Џ��n����ΟȀ^�]��(�[���gJ�S,l��8�=/�i�
)�{�:�M�[]�p�lq��x�h��՘ae�]q��#bE��K(�ooY	츕d!R�z�Wj������d��4�	�O(���l����	��
@��N"^���eg�p;��ค�u���B�B� c�.����H���KSp����$f���EA��*Z�O��ƈo�N0*i	|�O\:1p����T/��T;@��������r�L�AzB�.4��n����x�jm~��!���t�v�������'և����T�����c�|���v�o%��&��~�:}t��JR�g���o��즠�F�:��:YϼiX.�K$2l���of-�e{�v����0����_H���ýېm6P��^|� �\'�W;��h��S�<7̡$H{�3޼��i�S� �cJ��ͦt`��@Դ{�0c��6��<��� Dd ���Yy%Y���z,I�YH��*;a !�a������`?���{��)�b�����q�ɛB<�F��l~��8�?��5D6�9��d-����G���L�m@��?���K�g����6�C����h�?��M��~{���8X�N�����Mm�pf���u�c�Y'�pLCf$��-w�RJ�\�Y�[]�o��8�St�G����dz��Xgl l�I5$&� �q���;�r&��of8�A�F�8(���,.���	��}/_Hx�	��^x� ��+>� $�2��,�S>�
�����,�d��?�zj��u@�	_F'�!'`:�u�����~�Kb]o��E�7�u��?��c��*lq��F#!�����JH����4Q���1w�q`��>�3����[ Ϸ!O��0p�_�<B�[���c�\4O6b%#��҆)k}�i�Uwo(�
�% ŷ��P_],(���r�+Ϡ����dۂpf�9��%�D������6��9���&>�$���F�Q
�鉶&���/��a�be;�?�̚8}gT�Y�o/�%h�䗗���6[�?_0�+�����)��L"���E�<D[��6%�Ѫ$�sM�5�$}T5����}�M����g��4s{(��� OO��r�DOi%t�Pg�{.^�4��rn��E�!ƅmWM��[.١��?m�63����� �������;��/k��<�����
O�YR2&��gƴ�=����_U��t�w�x�ZYx�9��YR���j�M�(�-ZzP��{���`�q�aBXlxVHYEB    4f27     d40�2,��T�$�h	QϬ��Äu9����GYV�
�o�}�"��yf�k�KI�hWy�4����Z��<EO���ӭ�Q�n�pHP!Q�p1��k����_�����F]3k�9��'~��[e뜲�A�j�N.���mx΋ܡ��C|:~[t�E��bX��š���3����U�M�V�g�~����K��1a�\vʰn��FZ(|�C�D���'��M�	Ve�?��x!��zI�����7��1���_�J�6�i���%��2UwI�~e+��~�6��vۆJdwU3�r��/�Y���K� �<��1%��������S��d�2��r��*D���^N��p���a�A�
2�n������<V�K])���\���^�i��.Y0�#�D� Q%+�h�f�F"�Y��5E��-'�t��$�xTˉz��!90��o�dXi@�i����'B�����*h�����Q���EL�k�a���|�T�*����
�(k�ǆn�����b`?�����(�x��S�H��6oE�-!?&��f����D����̴��g�.�f!z
h,Q��i݅���A��0��	�dy2��f��[�v���d�yDz�ֶ���?@ ��hj����n���v����"�5�0t[T]����LG�TZ�^��i�����#C,�g6W��_WFН���d�Jt�n��:��Y��S��Y?h��n$"v�o�(a2�{�i�����)*ˤ���0V�N���٦�F�
�-�n9����*��1�3�Hp��[掉�c v+���; �������-BSU7�,��3�����7����+��w� ,R�������� � gBX3�배��}�˖��8�c�J@\����ũ��S��o��:ϓ�*;���w�����8���Ǧm�
�מ�z��m��yB�qª�@s�#�?��ٯ4����7��%I2dh���$u; �g���e�$��w�|P��8�L�0^pȵ��O�G����Z� p�.ǘ��,��	����.�qY[A�c��uKg�Tjr��2�~,��D��*�۹���'v���e��) I���D_�W�c�V���� �}E8��<�5wl$��+��߲��$�:����Hg�iϐ[�厌�_��{�F��	����ř�}�w�o����*gI:1�����+��E#t���OF������S�Z����р-
�'�!��ΩVA�.�(�7ܲ��5�M^l����gs	D/�ӌ����S%1��u������}� /��ˠ���A�sl a�Tiq��	��^���$&�碸:d[�@����Rm�l�DF�9LY��@"��E8�l��3���"Q�MRb+ی���׃&��PBs�}�[��~*���d+�6ICy�51#2m���a͂f{ײ�桌_m������|:��3}����c'�n��2��,��C��~6G}��e�����삠Wxvn)X�ӲB��m�z���*p��(�f���?}�Lc�?������;��w�ϾQ�z::�Ŗ1e�D(�p��<9��/֗��@���c���4���o�J���� y���'Sy'����ݏ7[���ɯB��c}a6Ao�~����y+c������m���Kb&G�Js��dF��W�@�Ǻ�ZO�dg��T�Ǔ�89���1���@�:)#�F�^E[��bj��PoX��6�cK3�=`�4�)V��sSG
����2�6��nF�nl�v��vGo)�/T���M���6��P����+���s�銹���l�~g42
�\�s$��/sTeZ��]Z��o9��b!URS�URް� ���u�9vh�+���S�3Mqc�u˱H���cB<0��$�|�c���m�<Ǘ��ДQ�L!4�$�=����'Y�N�her+���h�s��Б[1`x{�Cj���E��B|���t�cܯܹG�߲]��Tπ�2��x�=f��F�'���c�+�UڲHb�V\��-��������yL���̋�iF�|t�/�l'��x,��}R���g��m�\��M�3�X�N���i���v�?�S�r3IE��F�Q����{ Ntk��]w	�nм�|� *g���'[D\�e���8�"e�|<in��/�Ɔ�U����ڞ*�ZfC!Q~M���^���������\��B2*Dkk�QC -H�Y�0���UQ�>f�O8�}\Y��eJG��=om��h"���psz��@.�ߣ��杧�AG� �r�v\	���x��;��D�g1���z�v Y��bX� ��ɻ���A|�����Im)&�g�n��!��o/�M���u9�3�7��X�^� 	3&Z�֩p$���i�) R]u��Ob��u5�q=�����������*���i�����lr'����vpmb�I͏�_�	�{�������(�fɡ������z�,������VrK9������*��a�
ᘒ�U����ɧ�/�\_�Y�k��-օL髒W`���qR�-�?L��?v�/�Ȋ6YE�2�Ĕdl�F�eDٔ�޲O��6�H��2g<¥�*Y�6"��ǿoؠWD�{q�����}�/}��]��H����D�h�g �!&���.<��wNe&����l��	�ѵ�b����	\����[K0:p�6��`��̚B��f ���c��3�W]Ժ��)����#u�;E�i�@2;���)lX�7�������P_(\|@k�xY�#��/>��q��L=m��%_%���q7X�����#Q^Lv�g�\ͬ�pW΄�[��`�MUK��X�.�,S�Z%�E�'pЩ�E�u��[�0ܹ �MGTS G�#ϯ�C}e I��Ɏ6Ǟ���'��ѻn�R�j����(-!��ǌ�I�y_!ɣ�@�=6vl��(���.+��y'IH'G��0S��i	#&��`���==��䃄�H�ԕiU$e@�x�I�\	p7�av���=z>�/�yF�����%.5X�������"�R면K|!2�xX:����0��LnKK�"�Ĳ�]�84�b &MN�*�P��2�Q��;�.P�֚fH�dW��M��Z�[4��2o�p�k;�&8�Uv)ZyUC*�5�x�����BZ��f*H|zv>ȑ�$�K�-Z�lS�,�zNu�ƣ��p�gK	uu���j�ҼӚ��%���F����)K����0Fr���� {[��je�2��lO��?9T'�ާ�rAf:z��.����/���ӣ�@�-k#|}[{�i*,�t�o]%�9�bu	g%��+C�ϼ�R��FAzw�
T