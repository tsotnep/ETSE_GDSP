XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#TElG����F����I�����6�����k��v�73t�G܋+�Z8㬚�П�J�����1Y2qKrF�թ�Y��r������m�z
m�w�����%��w�H�4u��GfB�>� ��u��}�g�l�<s|�ʪ+:;v%��H]�,9{�MS� U��翱��D(�_�gٯ7�Mם�� �O�c��GY?؇D��;}��~����D!318��sng��-���J܃��A�e��a�$ \����dR�9SR�qB�MC�G��g�3�Ӭ�@퓆�!:��NJ!Ż�k�Wg�0��?=��:����x�t[[f�u�[<�(7�~l�Xf1l;�m"�FQ0K_�R���_H�Zuu��h܈#i��~���x3 ���ƴ��<��"�̩���d�f�l��{�"�����-d�fOl��X�E�q6O:�o�(7*�<N���A��_��M#f^��v��I��c��O2���a,�*N����.㡢�-��@��J�Ad�!�He��Z�lR ����.��x��\3�!|XzL�Itd��%�rH
	ț�`|;e
}��w�@�B�ʲ �PG��s7|�����i��:F������kl;���+1�1Q��%��FJ�aG|��Pf@�U����ݤ�m��zg���l��7D�����R�li3�.|\BF<��3oVD�Δ�8��#������g�����qm����ԟ�AG���w�:O=�����N����"F�>�l�؎ѷ��ʾ�XlxVHYEB    9de1    1670>��z��s�����F D�"�-���>�bR�Q���ѝ��Hs�7��b��N<6hC�P���>i8*��U��hƠ�J��i��o�U���	Q������m�s&���W,f�3��-�m�)���:�����İ��)�hA�66�f���(��-���D�Z�B�	?tz�ȸ0�����:<��i�O���E�c'�����E�[�o��������U%D{�B�/5ϙ������"����"���?�c�3��Q'��pԑ��;)d�f�5�����۷#:_��|���N���g�y�F�X4o��~�N�ś�e\9��y��RG��o��u�Ƭ�e�	� ����pm��aɹW�wޒ�J��W�S �.h=Z���d���lx�!#�z(��umw8������e9�B��=t���hX��j!��+�B�DG���f�A�����0mѲF�g��}}%�Ķ{�k�w�?@:](n3�Zv�!�(�m�օ~Fچ��7�4�8|��z{KC�*���s�@�j�./n��ރ*�CcrY�r�v ���6�m9~���6�j�J�6�����qa�Q���#8VH꿃I�a9m	=e�_����Z���b�;���^|�<���Y�]([pf�c��uU�+��/h�|��-Ly�	yT=?'��M����*�Z���\��ԝ>��߉ ����-LvT͵2va)~�=�d��
��f�����k��E�]c��V�Y��a�B�Mh�el�;-1�����%W��2��Sow�t���a��FXD&MAQN$�}V2ff�`#^I_��0��t=�7��t'G C��T���怓�����=����ȩ@�[Jd�x9�9W����Τ�k���Q8�^\B�tn�ww!����j��]*v`���-����Mp'�g��O:�&�k�N���S�L��i�;����B��lt�׿�sk8�
i��۹�3�y*3P��78��-�hKD5�}��m��+��j�25E�݂>�)f�:�Л<P��^}$]c����O��XC�lĔ\�J4����Ջ �Q�FP�E4OM#�>J��D	�IB��pG(���c$�r���ӭ�/�.8Ш�/���Y&,�1��x��}���_�Q�m�E�������,%�(e}�h`�$����J�}N$	�=Vzv�$�/m5[���n�����:J�+,h'@�n�|���U8&E�Q2X�����تD��L*p�&��o���Ǹ�wE>�{FU���6�eYx����A��j� ���MEM�HA�D�����>��i*8�<~�4l�����P�X������;6�lA�����Ǻ�����l�>b�t��D@� G�N|���T���ȕ0v��U����j��ߡn�Kz�`�Rev�}4�i>k�o����������_m^�_$��ǯ+ ��÷ݼw�h)K)8I%2�j>�"��"�$=�J(EFXv��=�*���_�>���#e_C�tvTR�R�dLB�c��It~qx9n�P�qu��vӌ�۳�rj�f��C��yI����0�@�n�խ�`u�������G�pж��NP�"���+��R/N�C�aX�@A��wps�{4Z�5]��3��<r>�s{�!ȥ��=w,sB�1�t$1��C7$��'�!��z���P*O�����FQ �5c�f3><�9���������<VJ65�h�!o��zd��>�*q�Y�ӤtB	���G2dS�G��%����1��ג��6`=��U�濾���&M-���a���,��L���T6M� �H��5����p�9Q�o�wYu�����
����9U��i�~ց��*�a�%��s,�=W�7���~�E}?�>1@3bV;V�\N�3 Eh�Ɯ$9w����cB|Laaj'|�K�;yF"��y&�E못��F3�0_�e'vTv3\�;�U�q�J[my�]21��X$C��(�
���C"�K*����_��v1/Q�"��|�j���
���#�阾�h�ت�2"�o}�Ř<���Z0fK6a���cow�7��`�J�Y"����#A�ɋ�'���|�F��i��w^�~�]j�h�����Ƞ(��� :���+�8�)��t`uiJv��O�Q7���;�Ǌ!�O��Z��{j��y}��t9KI�{e���C̴%��#]�i������<~��iz���;^~�g�4��A��%>�ǧ�' r)�Q4���_�V
�8�{M<�&}د_t؀���b�L�����E$z� fI/ pɖ�{�Wn$����Րo��8�!�:X���j�.�/-�ߊx��>��K�Ax�DL!����$��{�7b=�RA��}ܔi�ꋌ���tӁ������AFvx�!1;�}���8o_nr��#N4��d���Y�,n�U�|�'C�^?k�6:6+6:�.4�����/�ܤnK�j��%rd[�>L������*��a�q,b�4�k���ճ���V���&H��oH"c���8$Z���'�S*N���s�TL�q7p���y-p���]rJ�5{>���U޶q��0�5ș���v�If��$���D4��b>�i����S�����T�ᓻ��*�zF�,�9�r�*rY�E��k��U�2D��}L��g�9�_����Y�JS?�r�!ˡ{E��ld|9~�ݔ�G�^��%��h�����٥m�4F}��;����>���IlyM�̡�q_��/�0��?�?ZB��n�x̹π�X�!Z]]��S�>�:5��"����2MX�z �8�q����R�G��a|�K|���*b|�`��N��G�$x���"��\,$O���bW�Al�bX�\�	�o��>e�l���2��E�NG�]�����E8���|��y�/�t�{��FeVe��ogk��X=��̞z=Ӷ����׮�G������[ߥ�ё��E`x�����]��X�A5e.8�{�`����yX����V97�dA?�=�l��9z��#�g�\w\|�AZ���Q��������;d�"J��F�%~�h}�ܼB+��N���.�$�^N*����%%����  ��9ո9p��bz�:|�a!�wN#pR?M�����7~���%�����?����Qu\��A��Ss�sײ����yH�۲��[��g����c��8��������a��u@%����%���wN�{� 煈��h�W"�L�Y轼j�u^P,CiUI���]�O�p��>a�g����]^ш	D�]� :�ڞ��`*��`d>��q`��ڱ��z�j��qܳ���<�Ψ��'�0K���W�N�=r�2"�p���t��G��L�i�
�A;��t]압-���!��5�$�8TO.����ƨ��٩�ϔ�X�p��1E1i�����wR�V�;�@p���� z�Ȇg��
�yn����"�ž���l/Fl�ɼ��&���#��6�)�R��\o���E/gX@x��5���Ew����h�>a���T+�oG����x҄�L�G�lM2�i+/TAݯ�^��ঘ����c�u�c�3[�fO-��/��o+`h��P���~�dr-��W���cq=m��a\{�*�����.%�Յ�1Բ`H�������gC����!��f�˶�8�z?:N�0J�>�͆ܩ�@ٿ+ܰ��j��.g�|��V|�2� B� 0��l���'Q|Av����a��9�N{p��\f
9|��|f�����
�'�ny��� �ۆ�!��v{��,���B�[�U�%�S1��^����P����^�%%
��9��Jac�3NX��A�ޠ��(Q���la�C�Ʌn%�`F���ђ9�QN��P�����a�UGa���U�
ᖊ3Y���Qw�%<�z��1I��%�߳0x2bM�{Y���s�޳�B+{���Q�d��y���i#]H|��c+��0�������X뵏,p�;�uk��m��lP�����儚��W6��:�B�D��5S:��(�g3��f �Q;HL	�Sg%C��U���%i��a@7���|^$��Y����x�r���7���xL �w:�EM�䢍�N�(�-�od3��������|�"�`�=$�	Ά��Aj����d�J'm~�}[�¸�^��/�W"��H/� پUm�B�zS��p@/�%a03���)��� �~�ve���L�PN��WݠKw׏>D�9B){޵���L~��&Q�o��9K�ϼ��P%Z7�4]��!��c���{���ji O���DE0
}NK<Z\��^a�l_�^2��������n��\��@Ѕr=9H�e#1���N�yiڇrO��Yf ��I�c� �(�ȳ�q@4���"L�pj?Q{���#���f~�hה�ߕ"��_�j9�;u1�a��<g&�EV< �x�rȳ���hY��{�DT�8�ܬ��w�<��>��� N�/b{��o��.��f7��AQyn���j���=Õ����ݸ�8B'��}ZC�������&(�`e]�ǩe�	p���-�oo��$zS4FXg���U���-��1ē:�����z)&����z\�?C� 4�N�v���;�ĥ���F�O��R1��w�.���{���z����pχF��G(/��jF_L��r��|�������|�o9\�����Tj�P�:y�=͹�RGn����{H*1��U��2M�~6�!+��r?Q�(��1��x21v@1X!�O�9A5ӊ`n�{����@q �1Y��a?��+t�p�߸�M��/,$GȽbW���1��*Y/�E�r�}��7�NZi&{MO76�h��埥�Ci&Eo���4�q��%9+���A����`�:𰧉�+)b?�Ai�6�:iK�F����8��+4���|d  �0��#S�ysw4��?p��m�j`-H��u���e�I�˃�_��i�=�ߊL�ˍ
��2�M��x�3��"��v��� G����$d�QܑrNu��*�b�w�Y4I�_m#6����%�N�jaP	,��Kڅ�-��҄L���7l���[��\f��c�8R��f�>f64��G7P9o(o��G��ɫ�@ύ��Z��$fe���[��j'e!r,��3X]*!�
C�L�YѲ.�#"qH�J����Z*���vO��#�3� T��
������-�	���V����>�C
�iH�"�يED�R)�s � �����0�I�@Q��8��믒�K�B��LЂʟ��|3����.�\�������l#/-qN�7�����yF��m��ØQ�M�3���KF< ),����M���ֲ�ݧ����?�K���'�#�ڀ'�Д�x�¿8��3�_�����i@.�z�����Kl�������J�E�q�FIU�o��|���
��Z1�l��SS��b�C�̽ҭ�ҭX����瑄ϔb��G�iLN�`@��Z�&�^'���1ܭx�pX�����z3�F�\���Ɖ���Jz��'��ewWt�ޕ����|�z��i�t�%�J�c8Ȥq��"�ع1�U,,]�Ь���������QQx������R�l>�JA�JK�����3�i[[��[�J�(�2��5JPEEB�q