XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e�^id�?�j��%�	�!�sEQ�,;a,��=�A�0 +}���٭��I�2%�����~�8·�,��'��b��L95����g�l���+�3�T'4�,����(���4�����F�o:�MK����A[{���mh��zR�@���1��u3)l��Q�)��]��p��Xl���H(5N����YEQ??*r�pZ��V�,(0�6	���3u�N�U�Yї�t9�"��Z�V�a8��kA����z�P9�b�JeA�"������([��32%#����[�'JI�����z0�ԑK�3�lh$�|��ZC0����A�����a��|V�2=�[�I��̏ ]����GA���NT�c�B�N� �ǻ��r3�B���b%�^k�$��d�f�tDS����nƓ���T� ��E�����ߨϘF���(�0�v��f��=`b���|��{#�eV�u0H��`�kR�#.����J�Ǚ���=�e�xb�����»��丹��	Ҡ|�{�����e)ʩ5�Ge{ks��Ee}�3��i�P��JCUw��a�A3����a��*�=���Y@q�ka�����:�Vr�{U��uTŒ/|�!�HV�K�Q�	��?�T$=�KL��J2Y����
��?��Q�U��L����g���P:�����Xq�I5d�$�|z4Q.H�����!u'���y��A/ɐ5��N�-��,b S�{p ۊ��ƳNc�~�_E���)�I`f1���XlxVHYEB    fa00    2020w����2�n�H,vw�>�S?ݳ�C�ÊGM�\�*Iv�����~��G�o��ENfJ�(��Wx{� �%�D� .S��d�Ǵ����t�
/��S{��{e��\{>&�0 %�ag
���X� ���8= ��i��}�վ�n<��2߼<L89�V2���F��G��EY�4MI�Lk��z��e���VB��d3
���=,��
8g��x�s�k=����ܥ	3��#�X��-6����vl�g������Y�!��֛�V�D鹞����iC�Ob^_8?e�j�������%�Z(ݑ�(Epg��D���8h�f��& �ڐ)G垱���d�ǍTP_��ow��������������а�3
��
V���f��q��Z�S�ؒ Q�-K��O�)o����<�קV` YD�=	3�U)��� V�������/����i�L����$B	49�y�x"�'g*UHc N��e4�Ŋ�K���3U��zN����-���3y�6
@��Ob��wM���l��N��-�5�x��ȵs�iͶ)Y�$Q�q�����m�3����`>v�O�"|�[� �rC�WXw~1�+�W>�Hc^݃��դ310+X]��X��(/}.��@���&�pd��{�kD<iTx7 ���j�Ot^�U"l8{�(�;D<F��N@�p6���a ��Ze���B��i�g���99�)��Y�`��Nǁ@��L�
<�OY��*YYmDsZ �$^��
�G�'�,�ל?�j|L�,�E���֢x���0�6�~���˥nu��DoK��c�ad��������e�x#��W�a�x}�dT>1{K�{nރ�w�qI�����u�B�U��g���?�%�d��^C|2a �j�/|�cj��*�5��Z8,�7�.�:��-q��D�]���'���� ���(�B�٪��%��\M?]�9�JH-zk�m1�I����	�����Z|?ǶN���fJbD���^Ȫ��2i��o-�V���s���rr	?�_��C�	e����+�/�$7(	�b�P�$�pԮ�4�,�Zdt�ܺʏ����~ث�����]���73���r�Y��(�E�x�(�ܨ�[1Jڤ��K����cd�8�8ܜ�����49���m���/����q��j�����,�{+%�yȜI=��񄵯'nЫ������"˞�Ւ���/������6l�C�*��J�Q�,_ P����Ђ|��=$��'[ܩON�[c.~y��V2����r���٬�o	n��'���$2�Ĩ���?]������BQ�u�o�����sl�m��o���aM��Y��[���Ӡ#�DA#���3�P��Q\)�G�P#�ɧ/�5)�;D�O� �.�m�>m�&*��J� =���+7L�D��\t1yw��ff�nZʞ�R5��'"`�|͙-8�[L�<��$��c�t��W�,P��~�����\��W�V�g^t)��m�l��^Ϟ6U�Y!�{��F/O;7|�a.p6��������nc����Z%o�,�}���V�+��(�u!��?6V�1U��E���F/��賊�����>����Z�%X�#H����'J�I��� �mH�s��ۃ���i���q�^r⎡�j'�cUHYIu�6��@6p�$w��֌|rN���2σ2��[�I�+\<��n�p�n� ���3�����D��B��(��
,\��n}.���z�m
�|�+Pi�vO�^����pL�JX�綘!��kvjM,�����Wp�.���J�5�%>q�]-��j ��/�5�K�+޳/)C� �GH����ȣ���sWlYF��{��T/�:eYC�Q�L�Ɗ�mىQx�e�pG�H�=���Eߢ��,*f���R�?c�wu-&,�p����8��s@���� �H@R_���ٕ�(��������[#��6M8,II(V_&��%��~����V��
H���F"�hQ兴/I�Enyxؤ6�BJ;O��{�����:5��z(�F� ��Đ��H�쐋� w�A#�I�a�Rx|"O���j�˅t��p+�E��D��sag�G�Xc�Z���_<��]������\!qBt��VK�18ƕ��k�` n!PW+
�H{9m��7:/�H2�նR�s��A6,�b�e�����ͿG��V�ά|�n�N�����X("��n{�߄�� ٤}�a��#�k-�����7."\�6+�FE�X��KTu�߮�1�J�;�ƥ(c�('r=�!���Y�D���(#i�C�׮=Y\���m�+`��%����8/�:�d-��`عn�ƕ� �w/��2꣆�/j��c�se�Y����„Z̉5�-��S�
��`�ٴw����9�M#��nf��0��h�����(�������`K��\p/~f���
��ͮS/��Um����&s�7����?'^��V٘P~�M�P�K����
i�2
7>�KA�c���M��
���HnO@��ă5+��Ԋ����on���m��K�������.M���FrX<���d:e!|�!�}��j�g�E$���)�)�p�����s� N�X<:[;���ⓘM9��������k�X2+�^��m㿫L��U�q�Anf�)	_*�¢��E�;����y��ϙѷK1���ZeΙRK�������U|v�,�����U�X�t$�^u^�r�JN3|!U=5d�J�lW���n���G<2v�RXO�R�i��6^��n���b0��:ܾ�yX���a�*c'�(����-����KŢ`�f�ʖ�4j�wf�O��7G���9NQ�tkN8$�%��W[:�i0e�DR����t[q�i�BҊ��I��S$���mjB�BJ��؇�쮺���\�X�+>�GE��)X�a�~��6��s$z�	�I�fz���h�(Q�2���=�2J�!�>�A�3�;�GB�K����T��M��\#�<�s���C�#;�0�sB`���P�'g1���шW�I4H��UAM\�U��=�����)�����9�֜��O:/-��z�c��+O���ݼ��������k����C�k<]�g�3�nCgY�Ϗ��#)nُ�E��H��b���ҹ�#Ms��h�m�T>?&�Ga�	`�$ဲ�^�B�
B��\��� _��l��]�}w�s[�[Ajvoߘ_m�ζ@���z%���GS_q8��O��{�0*~�v�؄�!5-��2��je�0�<�<`��V�/}�l:�e������hR`[W����']�[��2�F��>��.{*ۗ��#w ��΄�啖F����Z��N@Y�"�f��:�g���IJ �";s��d7c�0�u�g4�4�{z��5�K���8[�]�~�f��6s�)��9�q��ǯ-q��c��Wa�Zx��"	�csm�5bi�b�C�
ߵ4BJ[�`���&�Ϟ���爚��T��^j�x;�b0�E+��t��ڌ~�.<=���D(�"�8"U<:��\���5p�;OU��=���+�̕1�+v���x؜����'����~�Vy�f4�-Li�?ſ�j�D�N�% ^0/`��VƠ�Vq�Pi�g���odV�X�0�I&��o{9�D(yZ�H:�0GgE�ݖ��6�X��ML��Z�����������/3���|	|�!ѝ����T4"hފ��Q�N���j=7jҮ�e
�Y͈ȉm̨2�E���T��y�7҂i���}*��0�k��� Z���$�t�lI���[i6M�|���ޝ3hiX�i0�丱LO5fP�V��ŵ���#\���A"���$� P��<|��7CV֔l�̚V��l/��L��b.�VB�*�)`h[�`Į;�6,	ꪙ��o&���j�MQ��%���閯C�6�f�X�V�/ы���߮}��ت���I��!�)n�1yMrb�^H��;t=�`�:k}��V�|uߛiX�\�㨞�⓪�%Ƅ��[�A2��l�n�`�:z��?��V�.�&h 3�k
���U�8��N1S�#����,�2�	�ēC�Ѷ.�Ń��i�ч1�7�R>�/1W�l
{�֝kߜ�!I	esS]�t-���mڟ=�����o,���ۀ��A��j�F*�E!�`�{ r��l�zX��L�_��@�S�b��w�.#*���'����4��a���Iƒ���GL"�u�qM�:z��z0��xw3䞅|Y���u_�N�>���Ff3I���@���";���"{����?�>v�6�{�l�}��o"#{�MϪ�;i-N�PZ�T�35X�s9��0�Fq�NtOg�ڄ��ީ4&&���h�]���ڮ��\<z�%&���˚�(�uq�g�̚�|�FL"�;D�L>!�D��\�yƨ8�\C9��>�fnce�MB��M!aiW_�Y�s�$[�x�݋�m����k�5�i��Kfq�VP���^`r�4��c��4{5�|��}�VG5���$_)񈦅�2ʗ��Kf]�B�ܔ��������	�]-c�g�*�J�"^�V7ۊJ]`MA��P?:TۄSyM4������η��$G��T��x�%�r�*�g��۪�H�4��4�7�4P� ���
q�J���'Ƙ^S٪��e+��ufMѶ��� �#ɛ3�b�����z�S�p��0�,��MQb�k QB�������{,����`�k6E��� ��C���m��h�B�}��� ��j�=��G�z!�_��p0����:XV�P%�m-P�&-U�J�����L�I� �����Q���nQb�#��e]�'���;�0w6���-V Qq��A��� ���L�/�1�s��Ǔ�h���?�����K%c�{��j놓^�mpQp��E�x�h��8��k�����P���;ԢQ����zϠ���7]殱��OE��?�lm�l3�G�b�C����Ly�����C(�C�G��Xol?
#ŏT�b��f�Di�.Դ�;�A�KsaC5-�E�fRG�bF���#_����h�U2���g��m۲�K?|`)�_R�P��2�*����S��R3�<=�E�&jٸ!_�fN�n�(?�§	}U8D}]��q��Ñ��`�5���i��^� �w(�Ѳ��m)i������5!�*j������TvF��w"��$����p�~�$5ײ'����
�����dh�j�L˄� |���ʪ�y��v�\�7�+�^��6m��[���\������������VZN<X�M��w@�/`2�A4S��~J�%�5
�N���Dx(���`]eh��-�����>�Lk� ��>�3v�(o��� �*Sг�u=�Ű
����e��%a����Ԡ��p�:	����u)UI���Q,�)Φӯ�Ib��L����*~v:c�(|�Y}�*�S�'������q܏�S���Ǧ����-L2c ��*�j�*{α�37t��{W�Z{�t=�L�jݝ�?�3Do�@k��5XS^?l��U�L��"�XV�!�W"�1�wpj��ʧ��'x���䔸`�?Z&�t�ݷˮ�`�=�����`��wg! '��L�0�Ju�ӝ�橃�!��$FH#ab�_]	P*8�7�ň���r���t�]9�ݾ�"���i����:����%VR�.�q�%�l'x�g,�� �mp��a⸁�w�Ӂ���U��ˡǦ�N�wE���@����򄩧M���p��B<�rx]I�Vǥ`)�2U��5G�ʰJ��<|?Pk��c8�'fI*�x��ٺ5yT�ǲrJ\٨�����-.���E�SQG�$�b���vI��p��C��F�G����{]�2
�Rj��C���y�ͅe]�N����Ʂ�{7}ĥa���9`���"Q���N��]�ɃKZ,l�pb�B2m=��H�6�+��kBٓ1���=AD���f�Em���/����j����S�2����	E��k���T_�}�}5� N��9'X��`�	K�����F���j� �jw�i������Y����΢�@��P[��[�K�u�����<L��~o.��&0czӷ���(5�Iq!��k�BS�>�'�,�W�l[R;9�_�ط�o�^�-2#4�יݶE�>�V�U-�%o�S���n0ˁ��'���L��+��'�uU��
Q�1xE��߽^�(���;��mB�g]]c�Ƹ���� p��	���K�p9���N�:n��ʁJX�WGC�f����,��֨�F�Oy��L/��
���w��C�>�����7���^s3�B�D���LJm�fZv��맿���W79{�B��l;#?OX�[>��p��8�����5}Fŋ;�3�2�ۄ̶ZK�@�#o�)8��X��I3B�չ�Q���.g����X�C�$o��t����ƍ�Tp��%84��d�+0p�p�����`�։nD��{yk�l������~�!!��ye_CdEV��!�;<�-��wXV��N�q=܋	��9Y�^\�?W8��~O$������ΰ�P8�#)��P��pp��@�t�����ƭxI���x�8=٭�uV�b��'U�O�?�KǱ&_� g��T�T�E1�@t�y�$���I�x��a
-͚`l�Y"�"��D�A�j����V�{��ti���yӠV�zf���}4���:���\�N��D�5Z�as t��F��������pnY�O�Q���H�v\��1OX����ƹ�=��/�gU�F�"S�·c��2�«�t)�/E$ƨ���CA�$�e��U�Hz��������q@��1��y���E�_���:6dl<j�7��ǖޢf� Q�/��!���U�Z��`s9K���]��VC uVa�����G=P��x��#3I[���2��\���"R#uV��&�T�%l�L��NPx/{� }��3�xc4L8������o��R��������y����JԘ�K	�e�.��u�S���_�e��eջ�'v�)Y!��D	�mXJ~�v����Ƕy�]�%\���� �^I�O�.�xv�	�Y�ß	��1���vB���c Pgˤ�֞B�H��)�[5'��W�6z9�# �1����W�:+X��}`O�� P��a�|�]k�����!_��Ϛ�i�Fz`��.��AkJ�����W.6����t�4�HAD�� F23�������L��- �EW�E����OS���-�;l�n��>�V�$)lm�$сno'~�pw/� �ޫ��9��ջ�N�w7��%�*o"p��~�����M��Z_p�H���I�	�I}�+/
�y �1lZh�A����G�nIX};%����s}*l�2J��PE
}��֢#�"|���N���5��Y�+z����;=p|X�镻)��K��r$���I��~�6i��@��;_�Z� p2��;�/8�>1�X'L!0O���6�灊 ���r���� I)�Ȩe���p-`�g93�$Si�˺��^���p=N���.��+�9��[!��,���?��!9:�˰�S���6�h�[b��OKC%Q9IcMVo�A>˥b�CJ���I�]���p�/Ctz��_�r��=vZW�����1�/Z	,��kxW�WkE����=O�u�/��9*߁��~����{��{�㶮~.�v	��3,����mӞ���7�b3��^��sy�[b(�D\�ۓ5G��&/$P&���M�;&��rБ��$��O$
P��n8q�潪]E:�<�ئ�JR�O�ZS�����);޲;������_��$ \���E��r�Q��=%󥣺�W�C�yA�ZMreܴ&�H�� u��:��L4���Y+	|[��5C2���!�/!/w�ً9K�+�~�\g�"�=�ʨ�Ph&�_zC�-��}F�v���k�>�P^<<��?	�&���0��\��f⟛��m��O��Oj��%܀%蹚�Э�鉍���%j𜙶�g��vtn�/����C�h30�8�|MJ9�?Q*�s�Z��!":��
V�O��tl'�N˳�`�f�ɽ+-Q�XlxVHYEB    cb82    12b0s��q�����V��y���(��@Ke*l&���э�w|PFU��å��a�����p��J]���7µn���q.#{:2H��)�h�������k�|�q�tI���^^�*�+�"�wQ�?�6&ȯ6��Rė�W�3[���ΫF%��ҽ��A��}֐�Q#��s�l7Q��Z3$��jZ��G��~��9 �}R��}����� 9!/���P��?�����Q��ֹ^�v �=�LTr$���9*!Z�g�ʀa���k%���6�嶑�?�5i��
�4��jQ9�z\���iB�
��"_�+���͎�s}�ಂ��ތ�d�$	?��z����0���{���$��-�����DH�9q0�0H�*�^�g>�JM��P��E�S��՚Q��&��C�ǌ�!oE�Z5�ͮU�"�"T�e���-P���C`��<,}���B0�*_�J�<���,�!����6+e:��yh<�\�
�d�(��E>��^{lye �ёx/�֬��7��3	����)����9��0	�Jc�]���3x��~��Ϡ�_0�� ��zF�^C��(��fh8�]�
��Ɣ2|F����^�6*����3����.�?���+�ӹ��;bBq�}��!&C�2G��/�&J�ʧ5:4����8�3_w?�pB��1�|��~����Ms�H1�ˇtE-���8]u���
��<�p� na�gȝ�J,/��j��Z�|� �z�8��/.9�}�I��07�v�@�^����s���;-Y�&Ĩ���Qs�ŀ��_,`�ͼ�B����Mu@��30��;zͶʕ,M�j�?��vٛ ���@��9��Z��"��Y&a���� ��ۗM.H���"��>U[����#U�����W1{��G����t)�;yS�������ss���$+����"��Gn�Y��UB�}I%�C_�"�!0ꂇz��W0q��GR�}!��ZUwe̿9���B<��z�+(&7�D\��%�"��uC#�cz����	Z��7Wy�����k�&8]�X��/��dr��9eޖ�Xg�����L
$S���. `��(�ؗ�Q�G
�<��פ������$��E��k,V1��#���x�%��p����qlo�M�Y.*l��Q�A�ե�i�Q�_Q%��wNX������aI���X���dV|� ����0�4��D3��'���OVD�%?� J�������:�� ���`�I���|X���{�f�>��;z����5�٘V(_����N2E�]�*Z��޹[���:[*���
�~)=F=@͎~hn�@�'S}f�#�տ0��Ŵm�A8�� ��~�ԕ�P
�_k�-�t��i�0�P�ZC4�޿L���g���^�v�	�E9��$�N��a$�̉M�����;�V�w4dn	�喔��K}zS�R���Au������%^Ђ�؄�X1�k_r��7�d0�Mpl��p"ڴ(kx��Ŵ��*&1�M N�&��oE��v���S���=����=&@��*��x�#��(h��Dq�]������^��&$�NZ�u�c)�9�t�<y�6��#�.������w���Bb?;�X�f��ĕ^ݫ3�yr���.$qs3|�
�<���F?J�k�wY��s��5K�����d��"�;-:)�h��R��N��	��0�9�eϯy�A����\�f��5������X#�{�eӾ���n��j���q\����,}�q��6Y�CUԜc�[vS�.���MP2V��)����)׬˸�����"��B3�2�� m73�gk��YY�ej.Κ�[�yB��w09�Z@���v]iM5s�j�R�W7L0�	k�(/2��Ơ�����0�P���m
�[YY+a�1�J�j-V�F����,��r��7���t�(���5�?n�n�FC�)j�=Zf����-6���&�ƻ�71U0W�6^����$���F!�r@�h�%��5m=g��7S�x� *�H�#W��yP���z2gm`��(�%��d+@�6�T9c.S{CV��!�$�/��(lO�]���1K:�+k/O���-�'h�H�jc9,ͺ�[���$<{�aHQ��l�h
$Ų�y���UqV���3�>۾��\��ׯ���l�4Hs�g�X0N�\T�/��%��Oۊ���?H��Rg�6�#���MG�:�6�Ư3����m�!���|?]�}�à��J�cߴd��2Sz�8��q�
�����<�p�xk+�Q��d��RZr'���1�0;i���`���R��D�q��=6ͽ �A,��Xع&J�l��*g0W��S�?G���F�i���N�63�DǁW���
9V�q$��Z�#�KT.j���2t}7��V����X�n*P︭��z �i�S�wޮ��)�$����R�a���5ș�N�QO�����	0��\��K��Eg�9�m�?8�k�(^�e;
���Z�{�Ȗ��Ark[�/�UeQ�$ןd$���'3)�h�g�\��7�8]W��
5������Z����T:<n�8�vU�zF��9���>Ĉ<@>�/��2c��z����N�������t�W�3~�u�稖�k��ʝ-�F�^���s��,�سK@9b���ӖE�V�!.1�]���K(K�/�)W����J@ב���.�>�E�L݃|���&y��c�/�s#�^�D��g�5<Gh�fN��r�J��aU����	U?��I�E���H
Yw�l���bB}���C��[�V������)H�m�F��:s���ʿ��7��H-��`�Yh�Y$C>�2�K �Ʊ�a?�]�n���Y2yot�Ȗ����f�a���s9_6���vr��BB��v!�RZ�u�Jg ��^l�uS�ѡ k>}�|�@˯D��ݪ�yw,\a�NW>���?��������>��~Z,�݈��w�t�H(���C�B� �9>	���4��d^����<p$�C� ���H�49�!|�m]E#��#;�2�����k��ZNLSv%�btܪ���&$m�l��N�����k�%J�0�N��'B@,�x��
-�;$�T�+�ϨK��w�$C?�}M�^��7��.��R�Ń�Q���KA@��\��mN���_G��/@vюd��e��K�[�qw�N}��b⨴��#�j�ϝ��tDT�R$z���	B�:��5��{^���8���x�ejx��A9")}ex�|��".>5nF�4���ގ�>���P��KϻV�a,�<a��K$�
00J�[u���\��HN��K��߷΃f-��#P �Kt�O�.-�6���T��y�I�Y�N�o%�o��k}T�������7�1'�aKz�T��!@x���"�ʐ��z�&���=����׍tw� U?�ň�!���&f�����Ixx�,���:����Eª��~��\(Hd��&�b�]�1Uee�Y�>�"`m�%_�bճ	��r�i���6��{�F/�#��^)�Sj�F+�+��zǸ��-+��`�L,�ex��T318��X��� ��Mh��|99�3h��cSߧ�67q�P#QŤO����)��RV	j�m2�/�s]����ևc[]���܅%3[��]J{!�Tg����.��$M�nYH�k�$s��:��v�R^׳�|��b�,}��T~!/g�N@��
�R��s�?�#����s���0��d��`�� 7���b��B�ԁ��f[�bp�s�<��2�[?n22����h��J�C���|b-u�,xK�&��ѽP�7F���lkП5��篕	+s��v��0,�F��u 1��h���Ji��ii(�;C��_:
�Ջ��_Z���/���@b��8��#F�[��U�%\�m���}E©�0��T[��6l;ںX	n�u������( *ը��1�Lp4e��Uv��栌��#�����i�|R�/�������oW<?����R�(
�|�/YS=�Ƌ��A��&����1Ɀ����v�_�����2S��_~�����}��-�ĕ�8����m�F���e�{�m�@� ��r #H�w}s��[;�I��J��<���i�������N��4�nH�L��0��6���-�e��f�2	��/�C��+��qo�D��Χ��ڇX���\5K�:�ѺOvQ�k)
k�w�si�q�c3���g���fY�ԑy$� �8��?Q�TW�.�J'����K�h��YiV��=Bm�o�r���7~G����P�A6<�������"���ǻ�Q��Y�f��V���� �Yz|�L��0� ���`�Ƶ|t�>��yR>��T�[����jo*n���x�v��ձh�T��Xg�����0'QmU٪P�Ʃ�U�'�Y7z�����!=Ay��'7�Dя�)���D��"䵑@��RJ��7��ň #>�:�{�7N��{ ��[[b�i)J�$��!vH�e��.��/3��'Z��$��S���a����,ۊ4���O��Q��w�cƴ�QX�����۶b��8��a����7j�k	6�-�*��!���/5c���38�{}�3��NEe�P�6c�&=��Va]c��}��	�6�e5�Hkf��À���!�B`��k�@+��ǀ	�wu��]���!I6���=�Z�M��S�8V���7�+擽 Դ!Ñ�Y