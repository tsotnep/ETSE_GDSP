XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����_\�$�mZs<
�%.�1-��*��GM�wb�_o��5����ES">[P�K'σ�����HӼ]�!IFB^��`��A��ƍ{�jm.��z'�?d��l�,��g^E����/�Џ͞-K�1e�cP�d!��]�K�~{H��k�ǧXp���ŘK�Yˌ�7�	Gf���#V��а�A������<������f��G���ɤxr��P<ô�_�S�}�*���C1~0���3<*���y�V*�(2*�\���4���D�P��;�ql�}�E����S܅���Z�:uJ6#]�mR,��E����� ��R��'rά�4XM�/�>��,k��s�Y=�_P.n��g55"����zE�i*�n��j|5�зQ(�����dY�ZW�B���-�:�T���_�;
�����1����g:$0��0��:�@�n��g����XX�O�~]��.�����r���X�x�;��tՓ�����]��W8��Wk�q��{A����]��Rm^��A��*�E���x��7�<FIcx����.Wl̨z�|�.mjz Y��>@��,�,������kZ�L@������~�mh&N��-�����,��yw���T�dG5�K4�4�C?�Az��:L��l��w{�����tm)�UV�B�3�_���.C�'���[^�E���o.~p����-��؍RR��HRL@�pE�<N1��6A�(�Do���C��؎�ҁ�?�b[���RI��EK3[�
_��'��XlxVHYEB    fa00    1790��;�'�އ�'�`}
��Ɗ�)�	0^���fw�.�� !�	�R�t��lQWX1/�ëF&�e�Tgr��]���e��_�8��=\��f5���TM��=�0ѝ�+��9e�{��-�@_傗��@���R����]���Db|�^ۙJ����=���xTY�5�C�K��Ҭh��\�����#F@|Ȱ��2�&�)�"OåfW;=����}�0�cM�eJ` X�b����o�=���?+�V2�I�5�rc���E��g�U���&y&���2���hLXƼ�{�{���P(���C�~I��"@q�;}��oHiC���F���;�翳|xo8֘'�s�Z�ר�b�4���K8:��a9���ݑ\c�r�pzP�g�y9	�Fp�~B��	�ypE}��U*]`��g�}Wkt^Tt�sW$�� ��M
"Q+�>�P��é�_2J4NU�lq��M���l/�T�~�����}��j��Ժ���SИ����p��9�Ҁ
+9#��(?5����եy�y�'�7Lv��Rg@F���:����kSJ�|��k��x�c�V������A�/ZMK�Kjž������c5#�n����ρ�\�����i�(&�O�0'Hzq���x"t�����������.�Ȗ��$ۋ�g����)�"���i�rL��U!=ڸ�c�'X�dg��ޣ��p��3 5\TP�~���ďd��`doRؚ����?*{�mm�����be8(k��2t�U����h��S���L�{�sy�]��O� s���-�v�9?���8V�I"�#�݆�ـ(t� $,�6u���ܷ	���$���d�<�lώm�l�]ۓ��|H�������E�bf^���QX�|E�3�檔hô�Ʒ`y�IK�ɔ�L�\G\��h�4o�;D��8��8�������5XC�ưv��Iq<?���B�ڮ���B	��E���d	�N�[u�SJQq�B �{!fz�?��=zMhnl)����O��J�,�0�#xy�������G7Y*?C�e;v	�#�a������`p@�E�M�]�F��s
��/��E��s���12tG����V\��q+�=ZGܐ��˗E�M҂��T�d�'Iq���fķ1T���>��q�3�K"K0\��7ką2�NT��(���|�6I� X�-�8�{U�@2J�0�f�z�7FQ(C ��VViȼO�S�:��WK���!��J����^�v1��}޶�c�E��z�s�BpձH�}1s�,>F*ւ�H�!+=DY4�<�đ�Ǽ�������HM@�r�/�?�(������8��wX"րq���N��v��,(Ȝ�t����gDB��a�Yܫ�������G�}X=􏽚ɮ�_�ו��TD�~�9ҍ�K��J�8�U��2C(�t�Zxm��b�����;�.ͮQ�% ��y��C����S��haqIvȌ�����}(�y�h����[��>�m��y<ݱqI����$]a�g���ȕI��uy~��yª�����`fI����1���H�Fn'K4���1�^c��J>�Z�d��	��+�M�_�ɥ̓R��8��_�q��B���{`p�C�Z��r#2E�Y�z���(7�����Bj&�l
�6(��d(��$@_��w~� �+=�≼ϜR�(�1eS`�$��%������Λ�(�5�$B�P�nz}r��=:@K8�Vkj���˾}"��I
̋Ea�U� �^p$Md���!+��@�*5F��$��v�\T}
���+-&�wk��U��ɔs�dd���b���%��R������ozذ�p�=�օY������I�G�U蚁�K���n$�ձ5�+���7K!��eOpV��D�@*SB�,#��(�S=�uC�C����s5�{�'�>��w`���Bw�h�Aw�������>[�����:������x؝˾����i���2Q��9S(M^����J�7AU�T�2�t�j��n�0�V&��P�?8�Q�][���~���{x��3�����F�~ )�KV ?��Q�ȭik��U�aug{b{����dC
�θ��;̶�A�Uk��@�S��p�h�cǾ��\^��CߺB�ou4��,�j���0�&���M�s�tBT��m�Y��v�����1p��Bom!�TY}!�=y*�䨰^̓�-b��a�	���d�1Ç,%��Qӯ�%@`Հ3������)�ˋ��U�%:GF���<�`'��*6�[�F�[��4�?�`��쇦 ԁ��Ě�Q[�L�W�0:H�)/�D/�7�9�����Sa�>�ǜ�ǹ�����JA��nz"b�4����3������xФ��;��8Juw�ygHs��5�R8\����~��`���s}�M�1�@�zsM`�:<��c���F�#mkv�ˑm�}0��)��3) >��hYE�q��tHGY��ٯC�E�Keay!�������#�\�����(�0<�%B0\��kgt���E"�!�?$�䀉�V�t=H�bl� e�������	�s��f7���cT��g�������׭9�&+�M��ݚP���՞	'��A�Y�������g�.Y�.:呅C�4��aC�yã֛�p\�cU�{�f%��(Z�~뒛傱vxyI�C�!�3s��3�� �̊�^����[����MZ�H4�I���ε/�U�\�����,b������w8T���m��4H��B�~�ن]i@��H�$�v��aSE���Rj�4'$����}</vȗ����}Dg���Vsf�dW$���f;Sd�d�6@.���p.;M��b���<�/�0��F�)}G0p,d U���b�?F�*�nv}��@��Q�m]Fs���{ ��S�Ȭ+InAV[fia|��|ғp�r1bv�t
�J��cuZa��pOD��c��� �e�0)Z�S����^&:�]������P�Io2��K�����oO<�&�|�\����w�<��rXL.��%�O���>"ۓ��L�;�k���Ѿ�gA'��R�.-�/�CD=��2��NF5ģ뢳R���n��8w�f����IC"ЌbHݟ�����%n���q�����y(`|B~BA$h�Ș�b�ilDU1�rͪ�h�)뻳��?���C+y��
������i����ٕ���ȉ�$��9��Ԁ>�U\�=�#85����a>�S�F�d`3}W�%�A-��M@�WӞݳ�*�O|V��J�ܳU!��
��Jw��Ssd�MܐlS�NR ���6�	�<���==n�$g��6�	�a�Kfby��-��Q�3�`nM�6���b�C��6.���w*p����	������U���e?��~�*���f��h�`��:S����sJC~�w^��4�RЀ����e��������-���$D�m�g=oH#�'�H�����H
�JWg$d[,�H�*B"�I@^|�HvI-и�0�%FF��A���b�^w�,:
t�?d�B�zь왊��e���[)n���TB��C	j3Mu%���"��V^����N��2uj��t�T��V���\�i���ڷg����J�,����ʗ��U��px� �I����w�}���//xe�u�G ���h �<�!�g��@9w�#̏Xj\+M
N�9����N_ݵQ�j]OZ���!�D�z�n�j4O��3�T]u0�J@��q[`�����sF�[�1��og@�6��H ��?���r8+�n����U�%-�]��!B����\B���s��|c�dD�)����ԯv��/y��M�zFo+�ˣ�!+ö/�AS���J���p��r��Z{� ,&#���R�_
&~�@E>�����ĝ�mW��V���@�	D���y����TýZw��ܟw��^�к��"k��"�Hڛ,�@*���L�ⵝ��py=����O�l��H��హ��<����,Dk���5�v^^� ~?CܸZ���eA�䰍~mȗ>�n�J�2��6�7���1a�x����41�+x����9mE^����2�bd����.�����Nh����@y�s/'{ ڃ?�>y��cq��V��F6��ł�ͬJ|����(�!�%�|NG�$𚴸HJs%վu~Q/������>��r�&o��
ܕ��~���������Y�D��M|��.�xfUF���qlcNn���{W�.X_��d;\�}�q �^X^��^q�U^��������#J 7%���5�Q^=E�����xL��y���DlȄ��d�!��F��LS�/{�q���%� ?��IH�]�0פѸm��d�lr���U����){П�c5��Ȇi��cG'�%������:�%�v�2	����@�0la����W��a�i���{��]!�����W
��K���h;�Xa��3�����A�Qġ@/x{ɒVl%
�R����ۉ�3!$���^Y#Tx"v�Q��Y����)�"(|�>�z��N��¹w���V�G+m�)����`�t?�v�JB���Y ���^	)k�j�U2��x���"����;J�dj��Q��¢�A�4m��9��o9�O&�_�4=�3i��(��ݿѺP�@t]¦��� ��Y��G#�
��������5���d_v�X���)�'O�㠀�6�9� ��Yʣ�\�ǦR�Y�Zn��E�-��sf'g*Xd��i�zC�`���6�������d���}�s�+�hF��v�����x.�H>!��k��'�S4�<㺶>X��Q[� +��6��ND���1���*���� !<�ͪe��h��h�b���v��8�~�� ��E�F�*�8Y��Mkñ2�i�^��dR=-�3qz�$�J\$��IY��,z0s��
�&�]^��X���������q�2%��*�-P����\b��A��sa���W)[.��ǈ{�04�b-�?|}	���T[w�KHM.���w�ek\(�����v�&���`���Y;tf���)f�X��,��$c�/-��;�����}wdSw��jI�UEBEK�;���mo�L��:�l�������?M�>,�cza�W�	�U�{X	��m�Y3{eQ-��g�E����,	)9$�=�Ĉ��Fc������V;B�tt�sk��L܄������Fk��3Λ�����ը�z�z�fxъO8�\���?�i�/S����f{Kz��A>��Kb�~~����� ~�'�7�[��x�ꂏ��}����J���r�"G��Ԥ<�����a�SV�(^�a��xu1�2��p3f�`��c�k8R�7�����PM��P�3��]�Q�D�5K��=�����d���o�X:<��ݽ`?��kq}���>|:�ꑞ�Œ��RO�׻$��{�S�i2�kq�.�ϥS-�;'�h���#ST���~<�tSK��x���ҵ������C:�g�����T�T�?V0�9-�ݶ�?j����[��Gf�ٔ�,�T�PB�P
�Β�7w���Y���Ջ�����/��a$ߠ�(z@����G�NFҋR �[���f<uE���)�t%��8ΐU&�����>���8�3��3���n�����̤��,82�7��U���O1�Ɨ��W��ּf>ys�[>�8A� �]�z�1��^I6�%�����$6=��E�:5N�l���4l�xM�]����ڵ�|��tE܃�fF����Yw�F�uC]���rw`�*L֠ŷ�H�	,S�R(\ڔ�'����_,p�g��$�0���g�xfƶ��6/�)c�mh8���Y9_P%q@^F>�gO��cå�Ikni�@�~�����i�����2o�;����XlxVHYEB    fa00     5d0\a�B�U$�MW��$�d�oҴ�h0�z26ϱ�o������J�P�
��F2,TA���֏��/�HG7T�_�(:�M0-�g�=i!y����5)�P�U�#�]��]V��ڲ`pP�[>.�L����҃A�Cg����Ke�$hE�DL�[����d́�(~䝏H���(؞`#T#��|��`ܢa^�tY�o������PE����A�Ix���uk��5�?_R�[�]�cqGE3�����,eJ���@D�2'I��S�ȳObs/p�%���q�~�Cv�M��o�*1��3g�)%Jwi� ���1��w)E����{�$=�%�3�����
f�!�.,	üh���-P'�2�~��oC���3&�FR��J1XWb�1�3詆&tT c����H�X������rf� ����
�=�h�>S�bk{������_��*f
.C-j&O܆���FWW��~�0�p/���[�m��vC��6�F�(D�&�J/v�Ѽ��#c��s9,/֋���i*��{�+���Z4�[��Ҡ��Ҡ@� s�����U���5xǺ�+���%�
��)��V�V��4*�}�����3e=zNv�jn�D߮�>^�j*�$�ڙ����[ú)�DQ�m��&��*kH7.s%�漆.����}�p\s�n
܃m4��С�RhFJ�@��5�T_5�"a�Pu���"0>(���-��]����t�ުT�ϝkx?/#(ՇH���Y?�M��Yl؜m��L*�ܨls�VE�Wu��@����1-6�s}D�fŎ�qᎆ-_>�s]�<N�~w��`��Ѭ��3���3Yg'I@���Y$��b ������]ж�F^W���M�:,B�/!6��W'7� �[d`W+�z�brj�i~�����S�#����F�?����� �Q�!�u�'﷛}:��%.n2��$��hh�WY���O�!��tjn	���	�B������J9	���FLp-����0�.u���v�L���`���ć�ʿ�q� �3�!F ��:�ؿ�m6+�P �/M���F$v�Um�v9 zz��uH���/UO�IG�&�:��+����)�wSAx3���Ygʵ�fD�#GvH�g�����)s�%�0�w��ouQ�`c�A�vscN�-ia$��C�l�'�"s�x���z}���rM
��Lm�9h�NwU�|������.�6�R"6��=����x���u�N���9�wK/�k�r�$72sw�8�c7�O<hA���'[��¨l����>>LM�-o������$���`��B8�0�G1s�(��~lڝZ�����(�r�u����ɿ�֒�f�H�s4St�\h�.t{A������q�N �4����j���Q�ր�3ڥ��P��Oſ�,���1n��>����ly0�����ݦ�=�`QοC�v�	XlxVHYEB    fa00     640<��h�a�3`�mu/�Y�2	��r�H��yPFu[�p�Np�t��bh��ψ�9��}�5�{�@��1)g3�UN����$2��;#;��J"Z͸ě�i���A����T�C�8{g9�o�U����	e�ӢV�єdJ�����LE�'������2��ѩe�Ǩ��.x�D�[��w�\x�wfHM��\Z��v�36F�.�H�n�U�(�����a��=�ښ�{���-��ȩ�&tTg���_qZ��7��~��㠠&�û�^�v�P�R�3�&��&A��[/@�;��gٯ���u��1�����4Z:Vr����,t�"���A���s�(���2�a'�̴�w�ȿ������4�6S��w����1�����{#�����^`��
�3�k��[)���t� ����.�R��!�i��[��Đ����<WD��YP��kr:�f*����-z"�S[�!g�]����7]�1=�E�48PW�;���� �d���e�5]�0I����s @g"%����N=��d���VKkg"��Bi��
z�GC�DQn��������b^����S3��s�c
�ް�Cp�,"Y�0�`�m�^��d�л���T�����-7+2���9����G�T���Y���6~���	�{�Dn>���`�s]aU�5g�~Y���D�7\��1�*��/�£�V�?�L�۠�;@�|��To�_���>��<�� ��)�n�����#���肣y�����\�6TɄ�Os��^$��Uq��T9MG��ÉW������F1�Ȑ�RG�<��Z�Q�:G�{jL`�ԁ6[͈dۙ�  �q�Wܜ�Ȯ�EĲ������5�51�0�7��f�s��v���Z�|��T��)(������g�W�M7C�����@"j�:�f�l%�ٸ���ʿ-��fH���bC����  �~��NJ-t��7��Iq*���p���9���_�)��f#hh�31f��_��8�N��p�`q�v���"zԝۺ^��/���H���%�0��� /�B���X��� �NQp�x����<��)��(�@���hh���9��6�'/b�i�kD#_��d;9ݾ|�~�WZ����C��\�[T��+eO�xT��q%b���Gb,K�}S�̽���ރ��-	d��������kJ,taI|8�*vC��(��2"�gjx�>H/�v�%�O�\ѷs� *MM��2��p���x7�i���'͖�'i�A/��1 �yX�|=�/�7���h�.hb�E2�w�t�_q/\�cvO"�&���&�3O�4�*�SeVoŁ��R��G�Z�&]@P���׋dg��S^2����LP.����% �w9�?*]��L�{���eAYjkb�l�D��dE��=�-yr|�Sq"�IZYK�b�^���,Z��(�Kz=L�����V�#=?�Џ�tܔp��H/�A�L�H��o8�g���obGM�*n��ˇi1%�v������Ai��X��#K ���㠼��[�,�m�XlxVHYEB    fa00     5c0�<�u��c|���O!�ȸ����i�$�]�0���DS@t�퓽:��璌�9+Jda>���x�w5���e����PA� �ϐ���ѫ��E��z���TҦ�T�n�D_��`ޒBЋ^�Q�MZo,u�P��ou!�;��F������}�)���K���2;���o;cϔpV����B¬�/�Y\Q��5j���_�7m�F� ����|,&�O�v?����a�l�IZGp�1u�qִ�A���,6�8�|߳���,O$����%QB`��J|�ݖ�?�}���z8��ϕ0���y�@m��2��fh,����o'�hP!\�4�C&����$��b5h\���uv�x<��K���Bµ^(>���e�����cS�I^�����4	6�[�Y��T�0>�:|��'X�!χ�����4x��TE�\<�02�o��64$b+U��x�@�g� 9���
ͣ�ph���_�$e��F�Hٶ��m�
���o�i��J���
����N�FJ�#X3P�L;ۂI�G��h���������T��1��|�wL5Ճ��� +�n���%#�P7#��:��u�"�/�HT��|��� ߸�k+Z:�o�4*v;�k0��׺����β�d �݂/�u%�Z��|�R�<���'*�7�Ы�r@ (q�rG�t�u��28º0Q����t�'>��xU�1����.���Q#������-�ƁC6�Rc1{ bZ�������Ԛ�h`��q��"ܶ�4C�n��By���K�׌�Z;X��Mʨ$#\�M��2ma�`��B\��V�i^I4�b凓ע����Ʌ��,G��}�KybOֽ�,����V�vP;���W�l����Ws��l�a����ho1^�G!��<��y�uI"��ԩ(#hd\�O�֮��r���f�������Y��$�E�v.�7]]�Y��2󯇦���b��WR������+dg���yʳ�7�P6Zޟ;��M�'��X��b�������?���,��D�����B5;�?��{�k���w<��T�^�&c�4��J��4C*N�;C�U�\ߨ;�͌ x�����:�oO�W:��J�bD7��p݅U�m����'Ei��&�f����=��+9A79֧R�1��b����sT�놹�T�����8���?�c��M�T����y� O[�K������i\U���g�qn��D��S0R������P'N�@��Sq��Y2Y�?�}�{:��}�� Ҭ!���h9W��E��p��Ax~�m�ưs��>\2��A���8�q�g�wK<m0�_�tMӺ#+i�,Io��p��w��a�N+���:w <��zR���:����{�~[�/_=�=�ŚJԊ�M~O��p$R�-�O���-�����;f�:���Hx����K�/� &�n/�Z36y�秽
�5�!��X��0�(XlxVHYEB    d347     a90���ݜVt�5����Rw��/6M��@�A�����셟��&�}Q�06�¬o�5� �9�+��S�ԙ�A�!�6��m�����&,q��O2V���i��z T�i�m�ߐS�Mل��/�}:�6��֢�#�JdOF�n@�Ņ<��|��pي>��G�q�Ąhaw춲� ֣T�M�/nj���rT#r�Q?�ɓ�T�S7UQٔ]��WP�@~���V0��v�ntc�=\���؟j�-߸�$4,������G1F��������S3�x��/�A��D�v~��2�F?F�V��>X��%�}E���N �����\�D�$�E����������Z���Sw�4�1��P6�q#���;|k<�wt~|���=G��<|��=<X�'2�����K�/(��Y=�����i4�;�9�������M��@���[u@`�/��y�n��I`#uG[1O����y���0V��,���<T�����c��=^*1��=�V�䫈o��SZt���ֆ��-�0��������IǓ8�AJ����fq�����g���D�	xS�����R�y��Q(
�A�0W��A�O+���%�<o���	`e���yN��YK\dR�eaO6/�ɪe)�����M\v9��'��I��/�)�s��jח8~��N@RA'��]V�]_�>�&.~Tq�KY�Zj"���`��j�X����Ӛ��|s ����=ǒ?�PA��[q�l[���f�R�8H�t�~j[j�޻�&�D39F�������D��^=C} dnOn���Ow�)[��a�R��ў(�3
܌s�|�|�+�IՃڰ1H���������+��\@-� �Q�������/~�h�x��z�fӞ"�Wi
L��\����!s�}�?A=)�(l�!��I�G����X�y&���§��P���5����RH(�2ܪZ[.����u���r��/i藄c����op6O�Џ�:J'���Q��n���aX%IX˸�H�c�7��-iP(��lEMx�U-ߙFNKV��3������g�Y%Ap�p�b\�����#��S�Y�@�X�#��1�p���Qf��QցU�I��U��+f�:��:{Y�V��38�)���^rS)e���HxbXҙ|ہ�A=S�+��#LN���y�ـ�ܞxQ���ٱ@|+�7d���� y�ܙ�Dgӿ�I6?��� 66�-a�[���9����4j��c�~0���ᬲ�|�A�\{�]?�;w�%O��N��j��;ߣ4��6pYLɚ6�Y3ՏHA�� S�N��(��[�
p�f��K���� y57i�¤�����j�!kY,��S�ѥ_�7����&)�po����/N�a�N�YP�^Mt������:}2H4B��L�bш�x2(1C�UЛ,pV�Ld�]R�>~T�ʪ�5/Wd����Զk�G��MV�TĿ��"t�q�)J�dO"<D�e�ס�x�B�f�;/ĩ��~Y;�%G��n:ی�h�K��ֽP����)��5`d�~�ԁ�/>��
�V����7.lSꛅ�.�����
�g��L�,��*����S4\�ؾ�+N��ܝb(����{�L ��n,^�nb�V^������8i��)��n�|�`�&gǉ�Q�Q3�i]���3�٬�m�Z�!,�2���7��{��F ~v���3~gA�6����8���pi�8bLlVm�7���W�KM�\Uq]P��\���S�W@R��.�'g!R)7�+��p'4w�\���CL8�
(A��.h�q�5�ܬ&�b��BZlx��Xw�l����k神L32�J�-�c����.�I�62}���G�j�����W�<�m�bZw��_�oi����ّ�]�� ~�z2�1����j��Î'%�L���^.�g��S��¨E�Z%�g��b��t�k%���f���p45ّ8�E�RS��b�V��]�Iq��e�������'�( e�;$�GXK5q%�~�^��烧�}�D�dAņ,@��
Ʀd�CiC��;R^����)�(^��2�- 7+���'����Z>�D>�>X~Z�=�&�^G��q^���D(�"��t%2*���͖��+���h����n�p�O�GŢ� �ygi7�����{��y���ѱ(4��z2	O���Y@t�+/T(��%�-�D�c�`�0�y�����y��	��>�H���Y76�*%�+���Q%?k
�14ص�7�^&�����cmѸ��l����΁x2�}���:]IDXo�T:C��%~i�����@�e!����M\�\ׅ�g>rqwy�F�L|�g��=�J=�Q�y�O��B㋨�b��,8�$ߧ�ʴ��Csv�&KN�2Ԁ�L�g\��m�eV���[T�CO��~-�=�>j`v�G=΂�ʾ�����Ǝ�#����йړ Zp�_#�l�YѠ�.�����QՎ�/�m�Hp�S��5����ê��'����58Һ�DrUX&�x�#���u3�YT �L�#������/%A�Em�~
������+��տy���?��I����m��o�}��}���)O�N�m�cj���+o��g��ɰX�@����U�)�H��ʅ��cQ㻽*P��x&�V
N��