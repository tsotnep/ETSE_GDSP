XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����g��h�[�n��P*�za�F!�WJ�Ī�%����EQ.�޸��G�>��0p�jo�.�{_:X}�Ӌ/��[Ҕ��%;T�k�"ЩA�]�٠�����/*Ѕͷߧ�K�5���@����*Y�E�y��+�
a�^]�`�o�I�����!�&?���:p���}�+;_8X�p��\ڗ��4B���x`�ٓ�L�3ab)���C�zɣ:Ϛ���1��7j�����#%Y�]�v�(_e0+��}a���S�Uٹv�g�C�V�c~uv�K��-ZRVl���k��n�nXF���0�{�~L|i�g/ɝR7R7�����Iҷ ����W�am���8�X�i�V��^�eU����ƽW���!�$���.�H�� &ս������2&&&�X�ۍ�`�uN��3N�2�G��b $�� �p&ZFZ�j�C�i��R��O�s>��d��L��I����/���Sf�Dj����/j)VV[���~o5�V�E˲���!�1����o����O��UW�g���F��7�h�t{'\�f�jYg}���']	p^�7��4��/zp��y
�W�kK%�ѵ�<u����!�6��t:��H�7 v���}uL:�"_�u��+��Z�jvn4�w=��Ih�z3����)@@�X�P_Z8f�pH7dt�[��,�w�:D�v]�;0��ˢ���{ᣲ2�`�<7/� �)$}����) ����(�����L�{����_������XlxVHYEB    9732    14d0�T�!Y��.��V�s���wP$���X�f̶��H�G* �"�����0��@�(	������\Ī��qu"z_)`-ًTy�"����h'���������:ė$�س�ћV�Z��]�p��H7��b��TUc�Zeͼ�JA�CWw�0�g�Kz3�Z����8��%���/da���J�k+D|Z���j]�葻�����d�l���SƊ��2ŗ.�=�/I�AU�^F�Ǆv/�N|RpB�(Q钲�Y��l�ػ�/��bZo������[zD^�׆��.���>�$�Z�:��(�����VO�]�����n���`L4��fy���P�d�F��nS�M$��`d�!R�Y.��� ��O��a�hWB>j�5c���r��w/@�̈́�{�4���*̪��$ȳ��>�S!�˰�5Q뱯u8�0P���`���w[f��q��B��bj�����z{N���ӵPmQS����Zuw��a��l�Gt����o�zl糓݀TkՕ�.ei0���of�v?�̶�4���&D,N� �1�p8PF*4N�Mכ,���%9�*���;�tݞ`B������5���uP��d~=? �;5^���Y8[k������?�Be��18<�א��x��I;p:ȋ԰=�8r��W��H���Fd����w�ߣ���Al'�:GO�Qlx8�9��6\1�`)���M���'%Ȇ���X��4 �9����:�%�Hb�$��!Mq�W0�/n���e�2R-��:��T7gd���y���z����E�' ��M��%7�����4�i�ܲ�%�s���篽zʷ����
ǀ�&���b��l��_���q%x+,�K}�a���N�}�ĸ����B��J�r:�S\܍�*#�_�?�D�ic:S�U����k����X�*y=���5����פ�uKa�a�F�� ;�W���8�I�j�(n��BԄ�,Ő�3�m�L��ҿ���
A,JB@.M����9 �>���ڊ���a�6�mBԺ��ֹ�4Y�{S������P�v9p�t��MZ�A�406��a��u��J��������t���o��qvloQز�gͼ�~�����܃T5�����C�ro2�ؼP�OhQCT�U�����I�g�*:q�ȓj�82f-$�g,���V�ߗ{VXFT�-�r%:Ps��Ɂ���FO�Y"���Z~����i�V�h�P`�D�$,��7M�a+����-�8�t�Xf��6x��XF~�@l�F����LJ���6J���~����R�A5	e!���1c��m�Z�^��J+4���m�\���ř��r4�MK����dļh6�_Ÿ�vy���v0����d��x<x�P���<�v��^��2ifv y�9�bh2��OL��~����ٜ�#ԫ����k�G�-ں���~t_��I�p���|�؏���}P�A�UFԸ�J;��M���/��C}�}�O�'�|����!T�^k�f����I����ʅ���Q-��\�&K5w�r;/z[8��ݤR8�Nn�wTY��^�����_�O6�UP����v�l�#q�Y�JI�V����&�tˣ�Nfj~b �)���l����v�(���S`c�qd�����$���J��2���,��)�Ey�pEá����kְW%$v�3dI���Xb��K�;-k�m���5��E+��sg%ҷyZ�Һ�>�6����S�n���=I�oY����>ˮ6�7c"N�Y����U6�\��o.U����z>59���	�\E�*��~&��L�w[��~��
L�����,s��|	��՜�gO'�
p4�8�(O�mi�m���� ����
7�Q�]����2�Ĝ���AJ��6�%Rb.�諳3%f�	�L�ю�f�H<���3(�$���G��DBؠ�5ߋ/�,Z���Z�$��L�������2L�	@"M걿���`���L�@�(0UJs��3��ښTl�	�`�yZ�ݨ$����G���� ݤITݨ�E��C�x�Z$�oW�R�0
�*��mll�H���cH�v���}��!�EdT���Inˤ�/J:*ei��*�6lE|�+X��G�R
Wʌ�w�;� �{����(a;�c��v��J٦j'3��ćx�J"41Ӊ��:�����#r,���*����{��`/m��-oA�:3{�v�#������R?�^|R����+��rNf@��
s2��Lp2�Y}�K����o�u�;��b�H#����b�a3��a�a�p͑S�oz�Q�EpͲ��+��a4l�M�d���?^���=e�C����W�_�{�w�J�����q���,�>���3O7�t�?�q̡ �{�HRFҁ��
��-ɸNB�!��;�g�iD�-	Sk�$s�#b6?'�����Z�E�'�:�Ϫ���[|Pn?u�j���^��@Å���a�l�t�?gPላ�c_�r$Ie��Ç�u���y����p��l`(����$�(w�݌2)�-5:��zb�F����q��p�g����'�� �{;4��8����ikׄ�,F�1��E���?�>"+�lB�W��� ߻�u?��6���4�ձ�&�PrQ�a���=QŮ�6�fԕ
�����E`Cu6��⬙=�(S��|ÿ&8nYi��X��p�YIi㜥��1%S�ǩ�b��!���r�;�_I9�#��(�
�%��{'
���@*
�����iOߒxQ����#�{˛_��	{�.��uiԫ�R��(l��ggy�
ז��;�7H؂�6��� ���w�u\?t#�i�����@�5ԯ��>��;����
J5n�6E�xK}хs�1ȵ�Y}
�H�7�`�o�0y�b(�Rg�n|�Ƥ�O�ل�,��	�i?��7=[�d*D�����4���i�X�0��d�81��T�]�r��h�UW���2�T���%�E~tE�t��ô8��
.}�k#n�|p��x� �3D��d��6k�����R��=����>X�1��� }�Ɯɀ�Uo��yӀn�wQK��*Ra�ԫ�K�׆j#3��a��'ɴ*�ގC� L��S��a����Ţ��H	��qX� ����k~�d����ԧ9䴋=�N�e�����{���Ur@D����N3�����zU��&���/"���,�}����pz0�hr�ėm{n��x;p���*���S��(U��8�����,�	`�>���N��,��kD`����m�AEE�ȡ1#&��!�F��#���b"�����쭫��6멷c��ON��uĈ���My���"�ܺ|Rk$�1��������O�E��:N�FO��s|��'�uw,-.�-aof�ִ�M���T�J�T��Y��鵅�s�d�Y]ɽ��4���q��j|>��]��'ced	��V-٘�X�rY�;�����(�U/�ʾ��M"p͗�ʾ�.gO�S��)y���{���I�-X���aqy���5�uP���;7Y[������K�=RS�����$/�!˩ְ<t�=I�e�"cE2/d_\A�l����@T���[|�j��(����Y�A����*���e��L[�=D��I�o��X��|~�����k.�hH�M�~
�0��*�A�tW����c)�@ ��?� �OIf�GS����~둱t�k��<�P�~Zn	��U}�_s����[�MO�
|��J�U�B�<ԾP��DEc��Y>��9�3��}�������Y�?��3�@��yFx�gʋڑ�-@"a��Rc��%�gGB{l���!�~o-���ߜ��}���k�#��o$  �v�����c���,B�����N�V}��ԭ�|�����hY�0q[ω՜xfk+��D'��E
=��r(s����\}cݸ�;��H	�a 4eEː�"	��O��X_��kd橶�D�Boْ�����ԫ�B�D)���7���{gY�l!J�	�P��m�p�����Z�N%�wv�����`"�WI~^Ry�~�-�n�O�]m���?>;�3�1z���P�Eߺ��%�{n)�"˘� �CN���X��9���	�3���� �����^�G��Q�sxn��������Pj\iZ"�v���΁���G��V��Q	 7[�\z%��q��Y	��@��fa�[7��
��j��F"�|��S�,'�� ��a���I�3,����Y�OU���xoC�qc��J<����͙{�Yj� �1������}�(4	<:������m<���G|����USi�����Ge,�ՠyي�p������:ؤL��;<Cg�t�
��T���i�?ҿ;��F�E�%�ig3ݮv�4�(�$��ͤ�=C̯ �~t$�F�ű�Y��2��)�m�=�H�!增w�Y�O��?n���<_�J������Z.A���*��?�O��n� >���b)hԮ{%��$7L8hJ��#�%���H&k�8:#7z�TщUp���8I5߀�uh�p��N����1\�]��u:��opB�ρ���̕���
�b��x1��1H��C��`����t_�����釬R�=�/�Cr/�B�T&t\����������QN��2�ݢ3R.�_m���S�|	P��j2�"�Bx��d8�i ۖ��6���[.��F�$`T	L� �{�Gt��߂�&i�}E�2�$�c�~v3c�@���@�Ԋ�(��2lo�=)�n�����G���5<�s�!�{���,HX%I��@�/tȗu��\��SY1�#�s��MY���pu�T�!���3���C�D�T�19XӾ�y���Jɭ#��8�j�����S��fpH��MT�:�&�f���^pI՗��I� ��V��Ȝ�BnC?E�R�6u�R	���C��g���A$�&2v?�88�3^����x����e���I�a�X�ص���q#�6'�YC�ֳ�[x�'fNJ� �OpLQ�{�R��]�88����q�{6�πe�@�kDk�3�gL-:��3x��o(e�p�����h� s=�ѯ}l�Շ�Z�������Q=��*�I�_l���GC͹P,Ǟ{��s�a���X+����#���� �x�I1�L���n�d`K0Z�r+�>���*�R4��G7��Lt�p7�hW������˗HFV�f�c��_���U=�6T�Y߮�����U��dȖ3