XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���y�N�bP�^˾N�n�~! �H1&���-t�łE]��Dg/�0�������l�@9m7�pF�oq��l�h�S�W��8��,G�P�h)A�P���y�k�H�c�̟y'�ٶ0����!*�H��p{L�"��R�L�`1L��@K�UH.I+�ݳ�
e��5�xj	�1�p�8�M��<��|2y|�{�.l��h&4�tj�S�w�-yk�OT�U�V�UG�x�5�T�G�����J7&(sP����=K�3�6'd�*9$q��\ZG7<�'�
+�M蠧�K�\�ώU���R0�$����@��l_r�Jto̟t=���xC�g�����f�e%��|0�S�-��pi�	�d���=!?�ɋ���ɏP;.m��K}hu��ck� �9އ5��{NC�!*\�Tw����3L��0-â�'�g�&	��	��J�u��hP�3x����*3� ]��Kc�pn|�FhG5�Ey� J+q�!�l�9ՙo�N��S,��]�YXW�� g20�����4c�m�,�(B��Нo�%�oI�K��A����A�\�)�?s��f�Nt ��C�}.�����Ca� ���,��o�휰t���E�MUa�r�rE�2.����BA���+�_�`����s�U��d��qAmNS�*��vUd؀M{����[w�6�%'��,�J�����hh�i�c��2���d�I�X��
*�x��4t��B���an$��r���"��)e��V��;���Hj�{XlxVHYEB    c3e8    1d20�
�@O
����X�l!�{�'�!����	i��#��A~�օ��)h��,���L�h��r }Pov���qf�6C�X�n?8��1h���b�g���/ƪ(&�w�2��A��QXK ic=g�N��	|ɦ|~m��2C�� ��ꭜ���jv�z|�.7�#3�3	�k�����y��|0����a��N/�0ߖ�?�v	��J�w~����$�oR<�Q\����:;� �m�C�������5>8Z�`�u��td_l�Ľ]��]��[f-�S�CS�����Vek��
A8���S�k�ǋ���v�%W�8��{�/V���?�/j�K�kt
��,�[.��g�Q�ǝNW91�e���ƺ���9�@�1s,Ԩt�9��`vEhݻ���ǌ��>5��+� EX�kp2��;q�|80R3ɩ��G��,!�h�8�
�����C��C�BT�rڭC�Mr�����d5ґ�e�!DC\���I�[�n�r��n�m�q]�]z���9�	_�aSLr��-b��c�;XF��� _�^��.s+ɠ�5�$�J܋o��B��h�	Bv�VQ��'�����B2JT��|9G��hO��?�T�z �^^\'�9;���s��B��/�߄�V�|{�4"�?��2����$��n�qd��J)*j�47�v*�>��#f˨�����F��F3�����V(��<��	� �d5g}�YD�Ėa:3+�����CɝG���R
{��Z���C[mA=/���C>Ϭ>�T?�!��j��Rn�WK��H|��(5�reh��K�����pYl�ӿ\����
��t��"|��S^٥po@��ṭ� v<��E(p���K� ɫ�=%N�e"Up�8e�,~��DSN٩Y�����L�\�:6.��t���Q�NͲ'@+�����t\�3Uq#MHS�"���� %٣�[+`�d�Io�^+B�x"�U�;��'v��v��'0*#�~M�Ř�S�=En��M����i<�{`cTlT������n�%,�}�S�H���������k�j�V�Qi �x�\J%�?���qj[�MYm� ;�d%49sH� E0ifu x<�63�Ѱ$u�_���q���p#�_�Eb0E�7�i�53��z�ɊK��?�<X�����٬|����)�;f�h#��h)��y�d�*fSI�+��M?�3� @k�&�W÷�+��0���)��l8x|���w^ꀣ���o-k��O���Z��Z���*�Dk���ٹ�i�B+-��S1�0���>Y�������퓴��<���=W�uRT_�n���q��^�c.l�f����*ɂڀ_u�����zYٜ���(������n��tu
%����t|Ӧ�Y��i�rK�Hi��É�Z��7}S��W �`iwu"��3�������
����+gV�`�9�����(���#Múi8�9��~d0[��hwL��iG�"���<�y-�r�M��ڞ8%��H��8��ރ;<��t�车���F�g����7�O1j�.fU���X��V�~�q�t0�5�@L>��o�t�+^v�Z/Z��B���h0�u��!�p�\�)�pak^4?4��X�0���jg�������!�)Ѭ���ᛄ�}���TW��~�10��`�������f�T?R~�l��� ]�<GJ�G���LC��H���[\8���V.�C����$m�.͸�Hr�I��i���Ոrf���"ՙ�n~`�G���C{��R��h����.���6�u?RB����űf�y-�+����.���D�#���ꚩ�A.��/8��Y��$����7�[kWni�7H	+)E�����}���B�{G?@YP���6���>��N�IQ�-h�h�g,6��Bv����� z.�&�<���nI*	�E&�ő�7�$��Z4Ȩ}�C������@��l��OW��J���o;� �fC�Z:: ��j����_�L�EDz�F��]=�{��+f9�ݩ
t���#��������bH� δ0�U��׻�p�e�J۟����'����������?�þ=R��M#���Z�y�~����#�W�<>3�p}n�uu[f�A��;�|r~��ť��:��cc�������<���9y��v9�� oO���^+���{NI���2)6���?�V9�]�&AHr�'!� �=������)W.�h�򮩷gGA�S��r����{�dx1���bx�)T1���{�&	�c)zl�p�Պ��>�>:�<���~���d��Q�����a>� ��`p7e����v����_��E~~�K���^�TF�Q�
��]�kp~o4�K�t�&7�`a�&w�oh���W@2�xHİt u�_����Tŧ�������g|�X�vB�s<l�!��]1p�#��ն�#5�����I٭�o���4�^��T��
,+�g���P���[�ܰa��i��3J�c`9<��uG�����V���%�6�� !0�~Cf�3�*��_���A�^➬�>S;l��d����Ǜ�0��.&l���"����p�3�4�<��$���"�#�}���J�HC9�6���:a������XB��S8]ْ�S$�^Q��.Z.���0mj ���?�i�<�y�c�����[f`��r��zq����-dc&�
^�"��l$2#�f$q��s&W<�Ѝ<����t��IĮr�`�^����vg:Cl( z�x�l+x�	vZ�K<�,�\�W����祐��x�D�Xւ�j�-�٦V������C� �M���5[G����xki��mK�u}�o��3��2|50Б�
�]H��e�/]�t��k28�mnӓ��-A��������e|퇇-�=��B���(,Λ�}�=�І/���0�=�e�~����m'-� �-^72.�s}�ղ���@�t^��Q��	��v>� ����ҷM��p��&p�9Ѵ��3W��-����d `��oQ��Tx�V`PH{$#�c�}]��2�p������E��y
(ebf��a���f�x������(����"���37��MM*sIG���1�^���N�*H�7ֻ�1�-��u6u`����#�K�|AÄ����`�p�I`s_�hZ��d]2|�Y/",[@�_
f9��)I�hgd�s�?`޷�ek ����<&�>Z+�kp�v����&Qz�%�i��ӆ������&Q�nV�Xŉ��Z��tX��٘�&4��%�-R��ٚU����?|�t�ߺ\�&W>8YGđݗh{9�}U<B!�z[q�����)���'i�Ҽ�Dΐ3jå1e8�ɏ��@\n8r�e2�@�G���}B�[/�>���!45�s�l���=��J;5�
��02�ިĈJ�߉���&��3w{x��-�]&m����rЍ��iM�%z�M]) 6�&���+�Ԁ�nb抳�3{�7OVy=�H�H�9��������7O���R����̞���yC9�\&x+dW�B�p�?\�I�h�MkAs8�| ��n����$�uʺ&�Ȱ��$m��	�x7E��m��AQxA��5Kswʘ����~�Fr�!χx]��6��F�u��6�\� -�>>Wq�Z�\���e� Z�����<`<Y�fT7����ah�_�)�5>ɖ�_�Hv��e��̻�D�Gx}��YPe��A4v;�� ;�z�;@o���;qTS���N^����V��SYh'�w#�c�AiD;�N�UHT�p�ʤ]�r���^C.cA��#���A6��>�<^�nTP�ruo�������r1��>U5�������)l,��ؐ~_����Ox_</8�2\�&�*r� 40�x�Aek����;��E$l��˼ȭ�Ù�k�ťSO�+U%<�pt���7�fʜY�FS����y�b|�9�4�$ј��h���ĖsR�wv����W!�̢�~-lkM2>���D@o�S� ��J�a��n�Hl��E�{���p;�s�^$�]�z��ΰ��0��M�Z-�|�7fG�B�q�i�j��לxG��FP��i`�o����{6�(�Yf��%����"�-�q�0���(*�%�w�=�/*/5��ucj/@�����Oƕ�1�����]1��H4j4e�W�/C���f�u���"�(|�S��Ǯ)��ݺ���qm:����r��]g������U7Y��.�:���
�����z��y�@��@��u�4'g5}�������U�Q�0shkiD��ʅ��q��1��\�d�C20�=��y�L�LX֝����wj�G�&&���(�P�px�S�n����'�� Cg��
�'�	�4.��:o���b�ki�8��S3Xً֩���鸋��X�s���,K�dK�J�%y9��d���4��8&��@czE*q,�Fxc|T��&�j���j�=5�y��o�4�l'�
y��ـoܠ��(�6\'(D��$;���-.G�y���� -&%��>h����i���|�cz�)�\�cT���>�����$|��^}n5�r�/�7y~$4?7U��Wc\_6�쬓j.&��xb�f$�8b6D��q�S����j�N�Lu�{���G�A�#y����ҕ�H�Y�x0����Ą�V1������*��B9��ъ �{z� ��F5g�<�ݣq�\�������sOu�(�?��,D��2q�5 ��]�J6[���_��Q��6g�٭.b�����I��ض-<����H����X3�v5�ac�����G߷(��x9�*OA�����hD{q����&�G�u��_����A]{��ڀ,b�R{�3Y�zqV"][[���3>��[�Q@�m����.�V��pj�%`��P�B���%�)�t��ѽ�E�o��`�D��d8�	���O�Ȁ��5�ݣ�8�- �1_��M���(��<�˭�������
�λf�p����E����72i��7��0y��&="�1���m��	75C$L^+�=�`�פ
z���_x��s�ʣ��$�b�t��Z�B1��U6Y,� �+������Ϲ�j>A(U?�F�%���ˉ����b*�*[�1�٨�rD*�M��.�6�������W+&c���F�B2�ĝ��JѰ]�k(3��)!�Dj[8m�Jpj�T��Vg�zät�vPo����m��.V��I��/{��ƫI��yd^6ؘ<R�ܦ�'�[��� ��MU#T����B�1���2O!��浼�9���O�
�t���W[p*hMW�H܈� e�ewI�ێ7��y2_�.��~��|�+�rs��qz�x���Ɏq�W�xL��j+D�I���pq��ӈ�
�)ʷ���y[cH��r03��g�*���J�8�U`yܹέ8�Ӯu/�$�����=Xx��G����Bu7�B� �y_�]� ߆����4U;L�t~������1�d�w�go�W�`������ǰn�PR�>���3B��>�4i`�ߌ�er���	-}�MO����<�zY*�=��Iߢ�D}�Pu==������z4��rϞ�Z�DI^Y�zХ-ȮC����ʡƇ�����#�v�r�����ê`��u�������˾�z���j�\s| 7D������2WZ�عI,�>��n�y���hj_\c\;p����ł`���FUIy���ې=�����7�D2�8�/�x�2^�o�#zw��������gY˪��{�wU��>�A�dD1܆�<���V°���gRc���'m��%�u��T�}��j�� 诐�2��,S�2�ȵ	K}[��ĝ��N�+��q8a�Qd� )�8y�S\��gzs��&�d�~��)����w���"���/��J�����?����c�P��P����mH���s2o�XGL�"b��	w�X�s�S|��AW���s������(7�fȓd��y�d��v���]��O\O?3�^X�L�f�S��!�|��;M� �,����QT�t�uF�S�3r��pٹ�G+�@�<�d��89)-x,���O�S�uыZ�BrM��&��Z���Gv��k���M���D��a��ʤ2+ʄ �:��j��%]$���rr���*��W��8����>����Е	\_��=�v���ĝ����ڎ�;�~�(п����lʢ����Äa�Y8�7������^,`K�_	u�Qx�� ��7&�#�"�r	���9Ƈ|soBVa�HY��J���a\��q�ix(x�}^���b�F&A�M�j*�f�C�Ͽ>R3�nC�2wo��T9��:t�ʛ��ܗ`�ڹD���Lr���ˣ�II ��:�Ⱥ�22�����2�b�2�׷��Nr�-��Bm �DΎ��S:��<_�~mK:�f*4D٘~��=/I��be9�L����������*,[J�Z��yIQ���� jj]X��3k��Z?`(~�O�/�zF��������ő	�॑&.Eן����cڿ��[�wƉ'	c[Z��z�~U��y!u O�)�1�ߣ�X�,����������E"�	�^a׍��nl]�
��w�>��\�~q�6$sY/lBK�:�{ ֘�������m�e�|]�n#�˧��n/�c��70���?�a䳳���fsiJu
��
6����qԇŠ����L?���Fu���&3EI����XI�g��`y�ْB��FI��U�:*:����	q �B1��!�S3������gWw5ʟ�`��W��	���!hU�K��
[�_��u�Dy����7f�'
���\HĪ`:)�ܵ���K���lq;6��"�Z'���
�c7�i�CL�rO��겔��A�#c�+��lr�H����t:��YT%J�Ȝ�T�ƞ��XY:`% >�z�{���P�"�DC�w��! F��]��I�$1 �]JL��L�Z�V��.nm,��P
�䐠T�X�R�P� �&�y��&k�Ǟ#!�{t�^S]2 $t��=�Ҷ�#��$ҔMd�U!,T��α��Z���P3
TZT>7��X��vb���y�F8M��U5�C��/3=�=�[���[�5t:��蠷����Hn��� J����������a'��E��$V:�_��M�hy���J���B���f�7�ߒX@cY���dX��ȡ����W��^�m{7������`�Z�5L0��$B���U��k����Q`�M�C�rd@G6|��,h>cE=�G����8;