XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u��&&��Ԙ8V�̱�/A3�/k��d�����`�/1��5>wG��Z�.�� �δy},-ݰ�n�4���xX�R��)t���AM����y{H�h����=%ށ�꨺@/�r"�^&����[0*��=rL��i�T��<("C2��X<�Q���k�?m��zNK�����S���פ��C�9��4���Jg�Ѣ˰V�_�b%�j�0�P/�A�����!EY&�Ak�kAj�V'w��{f��-Y7��;;�� �#���E��ߌ5�lgcC��7;xJ�qA����V����C9pO�z(�k1�#��Gs��F���G���K��1��r\^�^���wLF�~wm_H����v��5[I���
U"(�fq��(}S����R;.�
4}j�%)��B|�[�3�e�pVQ��i��q�T�!��2۞�(o�n���I!��N$���Č ��G%^�����D3�J�r3_A��;���C�u�:H����� Z��YG�0N�W�<�P��p��n�Y��,�Ĺ�_r�j��G�E(�)!.�Cf[|pr彍�m8�P
�Ӕ��`[(��{k�z��RX�-TzƋu���L�VJ՘����.3��a9��M�v��{�4���a!%at&�A����iQ/o������)\�@���^-OҴ
#ۻ�J����S����htD ٓZо)��6��p�*{w��@�*�Dq�[SM&	�Ƽ�#X �0��8��,��XlxVHYEB    7744    1780����w���W��'��y���QYWSNd��?ϐ���/��lgb�:%e�$��<��F{  RB�@G@t�@|��6���k�{�Jj���t̷KM�"��},*KBv��^FQ<�fi�l�wc�K�;�;�����i�'�B�d3M����10���M+ڱ��,( ~s4�+�?�|u�='9���&���v��Jx�?��۞ؑW�L��wm-��� 
#�:�e�Ӈ��V��ZP|��{f����xTy��a�ӧ��Q�pk�>����U��Ŧ�1*ѣ�?� �2KW��KyR�c�ؠS���	"�M�M�峉�~V�B�����n[e���  X��d��Owč��h���o1��&�'<�X���#�%lMԈ�G_ܼ{D�D`�Ei�5vo&I:?]���Y-�f��%�&�1�hl�FK�Sᳳ	��J�Q�a�����a��vEng��ɐ�S�����,p�N�8a���K���or�K��?�u�-�ȗzu
}�o�*˩��ZZ��2���o��#?r/!Bm��
K9J���u�4��i��B����4����#�%��h��}�#�k�#ik--R]�l]�+4n	���v����� |�4�dqL���r_'3U��8���=��op��$��$dm'�A����:�b淩#�g ������ʜ7�a�����P���2"
N.G��X��iw��<&I�E���+����m���+�����4/��G_���3��u)9���W@�g%Jpzd���g]"���yK�g��i������FD�}�VqB��\��]��S{��m�]4�8���c�V���OM_��ίS8�_�cN���oc_�9�=�����pcVw��ri�TP�k�#3ef(�{�F��h �>p�р��[��!�+�t��]��~:���X-#pǳW���HG<Y$[S��4����l��4}�b�M0"l{�	�ꉭ�|�		�g��aj�É&�߻���T�[���X��x�ԍ�AaЕHܾ�]��bT�<����yjrȍZWm�����x�8k2u���C,ˇ�Ti�13=���Χ��zD#.���K��b�+�<�[�>���h;] ����c:J)�����F�����Y��  b#�P����E_���z7�����/���?S�|��??���#k�9�l9}�&Q�M�񲮡c�Ϛ��u��CsXC�n�ӾOJ�߷6 �o�,y¥Y��	8]��qgWM�}*�h��_�%0�	�!y��_ؗ�*H�L"���g���E��͌��i8��"��HPɕ������9���Gi�h(W���_X�5��%��Zz TS�3����i����݅I�b�"l���`:��!C{�c���g.Ѯ��9�N��p�)�K��"�����5�_������݇C̅RLK��7���������� 9�ؚ�R�z�ݾl�˃6�flL�T�w;$��r�E��}�N�-��t(�����3�䞽[\��?�c�/E!E����.RP��p����
��k�!G�����zB�Nلٌ���L�U����/~��S����-h.W��,W��oC=�6�z{��;��	}���B��_S��z�֋댶]��a\nU�0��5��7}��@�7W�4b�ž2�JQ�����#����U�c;c|{�yJ<���L_Ө�!��J��_	�˩g$�y�N'��:����fn������Z�8�N�o8Ȼ%5Q���%B��e$�V��X�g�7�30�H6a��O>��-D6���A���Q<��A�u����x�"�&�d�(���uF[@��Zӫ�QW(uֲ,CF��mg�&�wa�E򐇔�e�Q=�f�����4>�y�����(�+.�yB�e�nиc������I� �������&�A��9EF1*A�� ���� �90�O�R',��q��D��N-J�x5���"�ȚZ�����J�T��6.߉��������y�-u^�%��耷��lL�jb3��P���1��q)�.xVp�7>w l�j�on�^�p޼�	E�g�!# ��V�ϓB�/�I�]u��)h�����(=�\qu�b;��o�Ba0��$����ه���\�wJ���(��L��x�c�X��O���~_\��#�9���Dr�� �-,N�ㆪ8|�a0����`��W�(����S��+&q�A"��zL=�j+���L�����f���C%�mM䪅S������d��ڹV	�xM/11�1\Խ��S�����':l���v�Eez/]�Z[��ߥ1ʆB화�b5�-/%��'%�0Ls����Gs����B����v�䜳1�%O4�˂6�z9s@�/gS�$��~�M�j�#����u��P�f�(�lD8����h�(7���J�����o�������!�;�~/��Ƴ���o��G������k@�N�$c<`n��ԈS��Y=Kz*���~p$Z�8ua����Z�x�>��B�*v0N7���T�@g�Y���v6��9� Hs�K�ؔ�?J/�nW;�z���=������^��a�u�
X����g~�AN�Z�v����.i�Bb��qZ�_��&=��~��s���� ��s�W�Gݎ'_JJ1S��6�M�X��Y]�F[��$R�:fP���4�;������ۻ���2?7��"�¤|t�S*@x�3��5Ud�0ghE�u����&��9��zG��c`�$��7���̔=�ч�y��=Q�9�k��G �Z��@�)i#\O�\Cr��� ��R���M��9c�߀	+U���KN��s��i��3���6� �U��aFO�[���������9��z9����@O1A?"}��#��^�����{h�պ�D�_��)�(M1X������v��鎄��|l�]`��ff��[��~j�[�>k0'�)<��QRt�D�U�T��ggS�+��[8FAO����w+ ���ϣ�b�����Wd���p�&-c�"�BPj�J�(>�w�_o8���Z�'�t�O�k<����a��x���Ŕw�z�_�n��x�����Ǫ+&W�_�]G�Ld'��w�����y=�LCR�:P�0���
�Ĩ:�:��/�gף��X�����1���*N����ӵ����P�㶼m;Z!��J���Ɵfg4im�dv:� ��~�w���Jh|r,�e�$x_����k@E|�Z}CP^c�F����V���¨�N� N@;�Ƈ�	�˷�;w~�#�놢�������\@�kVVhߓ\�K�H��Qs�A�ę���;�6n��r�B1�Yp
<\xs�$��������R���)~Bu/��A���@؂�0V.��U[ԇ�U[q�.|ka��2v2�G?����������>�Mn�T����Z�wh�fuy� 9 R����6��[-*�R:���k�4~Fz_5�Kq@��u��Q�XZ8�6��=��)Z�=�M%gd#�7\��x�l*U?�(W,������"��gݵ�K�;9��	��J�>u�נ0q���tr�>%�t2��W�H
y����	Y��\�gEQ����z�b{3��nt���z����άi_#��ť�&ɱ��}���RM�5i�ۯ��L�&�k��C"j��pi&�����ǀ��$Hv;��N����<�U}?��]�������#���q�(
-��2Js���%��pQg�`t�B�u����Əh��)A��΄�%"���T�2 
_w��o��Fu�����%:��y�a8�@��j��B�,�&2��[���{ �E׈��� �s�;�7������Ex�=��A���[ �����l����IG�8�����z�߯H0Df���uV��4�m�gh-�8;��N�]6�L{�)m�����G�X;3��3��q��������jnv޿ђ,���-��?��8�;9���]��������	�|�"��`��]G��>Ίr���YۿnH�޼�\��@�x|a����$+�=�k� �^Yr�Bh��[4��v���%��Y��v���e���C�{��X���&_po���'S�8��1'��$GYn�D���(�*b�	YD\Y�8�xf��wLD���� |N)��fD�_?D��G;Jy����%:rZ,��qY�
�����b ��~;K��a?/��|�}�E��!�E��󈓪�S�ʯ]�\�O�`��a��0H�������Z�)���M�T�bXb�y��ISw���U$�?�=��e�1�a DR�Vͩ�X����]4U�j	[QE��>�
 �7Y�MwTb�믋�������ߎI�[�簄3^��ҩ���v�DO��Q��y������?ܷJ������kNb)>��t�)���.x{ �
/q��]4�:���4�4����&���ƟA>v]G���ra�A���Ah `")�:-�b�IC9K�
�k����&�ɕ'������bv��Cez����a����7 y����t��ѥ�%x�@�;�4wq��(�Hi�r�5�)��N/�|�h�0���t��O6�⬖�l���x��IH��U�w��� sP3?o��c��`=Zu��/yS]���oxRY�&�����n����9��U�/. �<��!s`�*5�M����o��\OK� ��F�3lB�r?��a)�Q�fkD�<.�m�}�����r�R�[�KE�Lj=}���+
�OϺ;�o¤sLP�Da�\������o�����@�O#����\/�+�NВ��?�.tTI��P���T,�];�"$��΁�gIՅ���f����Z�H�8��-��Z�G2�fCVW�vJ@j7����}o�z�G�=im%�o�e��ʠ7��p��������d��c$9�PC&�kD�f@��E�3���ı��M;q��(|l鬠�Z��Q���}��8�]אz6s�q�BRY�E���~��b�ŧ�3ETP$�������_�]�Q�9�����kÃ9����w��*���<oWD~����V�d�s��>)�˒|�39T�"��.�T�/�p<�Z�)Ѯ�4���b��$<��K�.�թ\Y:��&nL/>�n�~o6Y�b��M�0��Ll��;Hv��#"v����x�wr�Q�Xx(�����^Lm���Lݬo�cVM��ű�>��IȨh�T�d��<�g��]�u���`s����%J���p������	� -5����6��:�\�*��,+��L��i��,lDk��� =�Q.�[�N�S����Y���x��/Rd?k;Ք�g��>�]g���r�l�F&\���1(C:G0g���Y��5R���P>�ͺ�fN��=�q��(̝�}Ocx=�G��#����'���H��>�4�8��m'�b�%����ѳ��vq���v4s�Oq����5�Y����".�Qmq�e�2_`������~1LA�[�:[ziv�gZفP?��4�����A�B�(��Q����Qk`8ɡ�_�1�}�F�#��s)YT��΢����?�e�y�o��y0��/�����A�M��(��lڰI�&��=-=A�s�k����o����~��ӛ{� R�Kf=��:y@ �&��'�u��=���[v��,�ƾ^��Cof�29�?�,[�E�q���Uf-kL(��Rq�I�7��u�ܻF协���h��_�.��	����kr��A��p0&8	q~�ۃ�h�	�FRF�*�	�(���H����Oww�>��� �Mȗ����R�n
$�o ܗq�
-Q�hw4WP�#>a�DG����} U+�Y��j8r��>'UW���n-�b�/����&�y*��,1�;���6k�z��Z������6�YL�b�̢�ɇ���>���ް{��P��N|ݲ