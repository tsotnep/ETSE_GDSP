XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�I��H�f�狮������9��;���FO�ycfʥ;���@��n��k�E����J͍����-����Վ�����|沱�h5�2�X/���C��~+�/J�G�X� 4NK�Q�C%�`�H�DR>��uB(L��O�����1r���+�e�ш��˗�����Jcu����lܴj��[�p����D��nl��9�Vl�=�m��g������ڎX�؅�ZY��3����$&+���I�q-���H嵾�6�������vᰎ1T6q_ e�'���7d�:t���(XG��^������=�'3��'P�'ߝ�r,q���^����A有q5{��z��v���!QС7Xr�0&^���|�VX����km������c;�i�Sѭ;0Ƃx�5Z�4�G�>h�చa�ް��U2H'��"@��u�ftϛp ����0�oEpS�J���=D�Ŷ^�&�kt�M���T���=:��H�/H��h�x�Pq����D77� �������d�۰�����`.��z~��H�|G5�85���l���d>�U*���۝j���͠���fM*K=>�Yt��5c���\����������xb�w`��0�̡*��Ej�����k5s�q�b���!>ڂ�������j�d�ڜ�w\)���DY��;DȠ�HMK���NOٛ�L��{B�x�7/��X6 �̄��s�<[�yH�*\L�%��}C��L	0�vY^�Y̲دk�� �q�XlxVHYEB    fa00    1fd0l8��NU��D��0����I0�$��r��ipk�+��-������|���S���`HJA�UJ���ca�aTiyoi��1��R�G����̸a���yk�]�*C�N����s��~�D�dF�ІC��=�5#�+���H�LЂ	~�g�Tg����G��7����%O:��Z���d5c
�����s<\|
��m��!͗@���[���	1�]1�n(���b�ƢRU������x���#춙Ǉ���*�׸v^����7����9�me�+ۅ�A��w�����-��q���G�� 5�����i�I���E��\؍#��m:x:���"���=R����-�moO�U�Z��t	'e3�9�膹
N�a��q>���a~��*u�rB�lg6#R7�������p�V��3%�Ԭm{��F٩g�8��9��47�`�/k�*��Hd����`=� g/��Qu���M&��_�	R<%'��`��6�3�g�`²������f;�:_��+���Գ� �һ�EK�AO.i!fD�3��������	FG(ыA[��M��»}wY�b�L���L�-��k�q&�rh�=��{�� �7�0!�[�|4S=������mE��c&?I?�"��"Fr��FpU6�l`aqZ���qs��X�����J��=#�Z��p���A4
�VC�Q�$�׉�n}+��;V���Z!2��U��rh(~�9�+7z��\fÙ�;+K
��p��_Y���H��R�F~?��PZ�g̪�m�{ʏ<ȶ)�b9�k���ޑ'9���J�9����M¦��*�,��g�T��p
�aVEn��e^��`th �Ֆ�j;;J�I���ݵ(X�]45S��=	�+y~��Q4'�o����g1���� ��t�eCS�u�����	������H�*��ґ]W�Vw��$\Q=h��%o�������K�Ǳ�\��΃�,���o����)r�������р���ʮ��`�j�La� =0�cD���3��ٯݰ�gʾ�!KZ�]S C���9�Xqֈ�.M}P7�e��6�1~��?������%�a�<?�*��t7�ċE�����"A� ��sЏ��(Q� Dʔ@a�(����(��1�B����xu�wg�Mh
����(��(;up���v�j�����i�w�G����&Ï��ۼ���Gd0�g��|�ڕ���S���FD3����n5H�Y��đ�J��?[������9G�Q���?��$&�|ۙIIO� ����q���������J�sG)���GzO�t��T�a9��x����'���R���q6�.}�}�Ot:�%���8��!�(售w�d� ���#��b�Yc�6.DT�i�W�ikq8�V�y��!��ݔ�<��x����h���e�q|�#�][V�Dn�o~�y�s�-�v��N's*/�LY��֒�/�oD�Q׺�3���B��pqT�?���G��:�E�'
�rO���p�V%!a��'W�z��4�;y[Y�������Ja��;+˾G�/���,�7C��<�sr�_�i�T����~��F}�3��\��N�Ow�2����m3�F�3�Ep��Df�8L�S__�0�k���y�Utd�dO� �S�4���:�:��G2P���(�^%%�aK���	���m��L^�F�>a�.'_��T/J�%�q�h�k�i�u��&�Y���%��e33�� #!�Vt��1�k
rZ|�8[����?�U��o��}.��Z���^�8mBr:��
�z]ݼjL���?�+��r,}���s��E�<��jڄ��6���EM���%��ǃYWR�RY9�7��Q���8Z�W�R	U�2!>��Y���~��$��x�0��,<�f@:�UT.�dp[ �hr��b?�*����*�5��,p�;+�WC�|�o�h��\��0��w�� -��*�ws׉��m��C�u��'���6��<0�٘�6��r'���ݰ-��6n��-e�[��a����玕=�q���I)����������:���rBB���D.�	�X���RKÞ�%:��gU����*�o����e���	�9k��/~(g .�H�9�����V��o�<wdj�k��S�A[-�i��$p��[�C_FCs&g?�Ǟ�h6Q�����rqh��᧝��sX����Q؋˛�0M�l1Ũ��lV�(|kq���TZ�p�a��B��^Ea�f���[�D�9�|Ȋ�gB�,f
d���u(�~��%|cH��p�;��'�i$�V��^�k�A����gAS�ͮ�ױ�U(j��:԰��9E��8"�!0T�_{�No-�~�b4{3�C����/c����U�Q��L�[vmJ}��H�Yآ�:(�m�W�n,sJ/剤��=��Ν�$�x�_N�m�
d�耍O��_m'�~����.m��J���_G����7�9��e��1��^��o"��6��^a8��,q�W��N����?#Dߢ�����܄��b��!K��,�-�vsI�F@:�}T�����kJa3ka+��]vE�s>�V����0���vVL���,Rhu@m�i�Yu�s�X�7 �t�J8��j����<b��U����/�I�颽��#[W�ى�h'oÉh��xl�7��M)�u�䔁h����5�U�]%�{���+��kn�*��Fdg��ؿ���TܷS rse�f����5ʤ�lM.����:W���*/�Q��4ɩ�D7/�2�����h;��z�/%���x�vF����F���@��ؓ�M=� �e��)I,-��@<����>E��0ؔ�|�O�<�W$a � �x�.BF�$����պ���Kj$�&SY�A�].�*��$��={؈r���9E��*~� �5sE��u�C�W�Fj��ނ�n������Ggʵ�D�	K�x).�c��ڋ�z�C�+�ّK�?�Da%���^_�Ya�К;-�s���=e�cU�-��򩁯"�������%U0�aC4���Oj�u�9���ő�j�A�0��� U��V��0B�프�|D�����M��W��K������=����d�.a�Rw�`���;F\�D�
�79�P0�T����|�6C�OpȪ�'�ȭ� �N��-y
>�D�Q�G��e{�By�g��?��� [�↵�X�E��=��>�fI�܅��:�o�PO}b�?��.tPJ�D���-��M�$��x�y|?�f�5�Ї�B�u˅����J��� ������#���r�,��Z��l��U�e"m�z�\."�Vq���x��?bqתX�����W���o�^�g��U��P�-�v�L}��/{�}�,l������^�K��8��Ѱ�&Wn�&U��)A�C��a]��;6��W�i�`Z�䥵O�:@���S���l+���X�Ǻ�33�|?�p�gkj��$�~Q1?����)�}~�8s��[��c}�h�W�� ��T���,��SC��w�6%E������a�cm����g{o]!�Z?T�[E8�1�����(f���_�[$���5��)z��#����[Fؑ��3ܥY(p&�eW�v�.@�q��2�,2Y�kDT�-��KW��l�7׭�ƞ*�I玐�����%Ѩ{nDe��a~��;�T7Ćc� ��Ū?ǀA?>�C��oc�}�|���Q�~��wڕ�R�u�N$��G�7�L��la�,[�x1{p�)<��HA��|7n�!,�������|N�@i�g��G^
�+�p�)�w�+�Q�'AJ�_�2�/���fWB >}}*�HW%܅�l[4���J�tQɿ�Ė��V/qeJ�٧Zчь㘗���E��t	��?Z�t��$�fm|VÈҁ���>���Y�t}Q�_u������a�qJj�Q��$��8?�FW�!DE�y!@�͵c�����ݮ������r�:��u��h]���f~_47ۃ���2|�����&Y�\��(�Z�v��}�[�"��Pu�vi�>�z�'K��G��ql3�1���%n?��3�u]�ǧ�q� C�
�6��:]i�<d#��߬����sm���-�f#T^�Ô��ޯ�	��é2���G��jyv��m,�T��X� �i.Iw��m�
�L-=�  !E0����݂-V�zQ&jk����^h����hR!@͑O��a�d�P�J��/��7����t�c�2ި;�(��մ�M���#�h�h�Xy��cGsh�U��R�x(�T�5��B)75LY�[���%�c���#BB-�w���f�LN6+Ւ���xpp�D��+����k~�>q~>W�1e:8&{�\�ܕ醷g�RUN��P{9ө�XA�� �����4nP� 
�����f��C��>	�9�癎�h?l���s�����ʻg�������9nlG���n5����s�'�ms#�L1�y�3T�[���'�K1����h��[�:�\�7n!f9�<pU�ٍ���'s���#�d���*<Mw%zwW��G<�ZQ��b8\`Πn̦l� }�.��&".t�'ID�;������x�~R�s�e��/,�G������a'�B%Ъ���=�6u$^�;c:��\�>=M�K):����⚑򼍻2ʡ8��2��f�c6�^]V=d��7R�ܝ9�aG��%Z�������h��(3"�\�B\1'����M�����rM���2j��* �� �J_��k�O��\`����ʬ��*yJ�G`���ix�ִFݝ��&��o���a��I�r��������[m��<�
�K$i�C�2��0?0>a�ϐ\�$X>�&`;�͔5�T��kH������G�Ӣ��莮�e�H�o��k��$�Ǫ��~�mU�HjmznV�0#I��2���
�vi=�@I����F�L��X������	c�ץ���x�H4����FS&�Xv�hH�Ԃ_�������:�j�r�Z[[�-�W�v�$P㉹��h�k��Aq�#a�)Y�2U�z���0�����s���$u���hz�s-���c��[aq�5�̜X:��C�f�Ʊ�l����梅���YX�����ݢ[)2��L-�٧�#�f��S�ͯ���B�J\�\Ũt�~�����5��c���2|�j0�S�ó�vw u�ݲ�3�Լ�紤f�㿯�!�tv)o��x	�61�@��7�)�d@ݐA�t����c�w ���̣������f�����&GX�Fr��KH�����>�&ڨ8�_xE�=[뤫��h���P8�慼��V�F�;��H�N��{+���j����,��J{^F0��tRcL�	���xrT�t�i�vƐ�N�yz4���6�,�*�Y�欔����x�+`gG���ߦ|4�c&�([��Hށđh �i�Ϣ�F�w�?:�i��k�ऻ�}x�$�_�$<�;"J��`�t���).���E�����<p��`�{c~#y��/v�W$�7-;!Kf��¯P��>8[���^�Y�q^��l�Ɨ�LXy�-�e�r�!H�Ћ�� r�!�i,.�d�~إ,��5�IW6)���y����.9E17�6�=οz���}�~���kt��NX�q�����G�T���i�p;�F�3�o��[���5�h��0�)q�>�c�#-� ��m���p�j�tZ�d-RXK������ߧ5lB�勞#� �sBs�����o�0�&��eN]�֎qab'4W��/@?�h����t�2���go��r�WH�}�]T�6$��,,^�����r+0��֌�颰-s����h�R��b5s���.� 3��h˥���W#)�y��p�ګ���䦫����"	��_֯�/�"�p�	*� }�\��e筨J�i� �XU���Oa�o�A���hq��g�Vp%$'@q��F���K�'o�Cv��𳝖]�BR��Ѿ�vq��A`�8ѭy+�ڤ-�A�ʞp��ʺY��j^(�e�8��{�8�{|��:�0�!�p?��/c0��dB-�����^r��,���Ѯ�ŵ5�vޥ�}�|TL��Τ Y��H��S�,����u��z�C��d=��Gc�E4�5{�̓o7ӷ�Q�7����b���]
�k%ܒ��Θ�V�A���煰���A����wit�I9Sฑ��V�0��]@���41G� �o����M�,�
]@������Y��E�Qv�կ#���J�#5�%�g��̒����H Ҟڏ�·�ZL��N�Z�<�`&�r�:{���ɩ6��:ca���z���w!�̌F�
5�mhJصB��~���)��J�1\[]<Q���rf�����2��%|
����ph�rn�/.7h�Q��H=6�\�F�$�v��(��z��&,�lmZ����*��m3�@�s���V�8/-�=S�htF�$5��b�<^���3俹GX�U�Hu�����d5�����^��!c5"WG&O눟P�pZ	|AII3���Yҟ������Iк�1�� ��&��@�۩r�<'� :I8��,�q����=��q@���nuL�]�0�y�i�nցX��%�@qdp�����>�)����������li�U���5�Zї��m��<��lK����qq(����h�@���^2'N�q���_:Ym�[��2(��g�b�3d���p�A�T�Bm�plö;�
x޿]~Th�Ԭݢ��OU�[����?�{k��E���O�6�?f3t-����$����{)��G�L�)��M���\b�8�B�_�H>v��l©ke��Q4o����'��)��@���M	�n$�$�PW�
O�2�u~meF�{)� D�n������u"_rFEm���ұA'��s"9I���^�v�����f���wA,�d�=T\�da7h��7T!�ҷ�L�}!a�m�����M���0uAñŇʃ�2R��c��,�Q��EŒ���)��`�.-��!���5*G$�a�i�
�N�D�<���Ղ�rSi��"E�u2��\���c���1������2�U�t}��ٚ4�p*O'��b��d��}O��E��͋1�E�N�^���G�^����/��Y����d��%���d�-y���DM� r&=aY�+��`�������
�ɚ�$hhT8�Ov��K�u��!�q";O��=��suq�$'>U��_&�D��� ,�v?�&�0C�6ucW��
y��K����5�-�n�B�S]
��������r�������$S�
�*�8&I̼�W#�	[��61��G���ְɞ{���5sM��尣�G?��=+ђ)�)�U���*`TGuP|"Qӵ�k�{fIH`�)�t,
�k9"jߏ4��	\|�!�t@"�L�?�:�Xpզس����ϕ����-��j�FJ��j72����[����i5��>A緊�U�ix���Q4N��%7'M~���@�/�Ѽ��o�OY]^��'���.s��oR�[<�o�i���ö�-Zh���x��ˀi��k����٩R���>��r�f��1�K���޻jt��l��5�f�a�ْP������*�ώ%�DߧK�^Õ�)�����D �O%�vx��d
#�K:d���8yb.�P�C�E��1�!)̕�A#E�q?5$L�Ԍ�����B��%9��$�]5rs%V�3��-��
��,*F�*-���������Y��ײ;���l���g!?�|�w[����3��bK���[�5`��1ϘRBMbf񴫒��]��K>a�;7���"���1^�d��2p�'����%!]�.
ޠC�!9��┵��V�j����;��B+��ʋ��sl>�O���ۡ�8a�VD�4�&�h�:9�����]��S��"<��Dp��H9ǧ�����T��p0,=+��i��U�j"XlxVHYEB    fa00    1340gȳoӢ�ܻ�r���.�@i��b�=fy��{VF��\WXdt�Y���$.�:�i�P�}\�e�z�ۤ�~ʾ[:���{�!�j��X���ɭj��F��v�i��/�1N�*��2�J�U	�]����	�G
- �ib}E�u�љ�C$���K@��/�|hk���ڠZ��9Oڼ��Y�%эFr�8��*u��*q��� ���t�ͳ�
LYͽ�l�~%���m�`#\�Ś9���з��<���}B��1�4"|S�we�H&����d�K���ܓ������@`�~�}�ڛ��&�����KͿy�i����<���յ?�i�s�j^}l���u 	�X��|�H���Љ,��=��f�;>i-}�8(M<���k�\�nhந��F��jj�ϼ�jC�h<���އ���y[�	�a[�UK)d�깤�K"���i���y�h.����
�^+'Z����}�C��ٍ��w�K~O<H�o�=eǵ��E&'G��*d�t"
z�V8�\�Oc#���۪?٭���&@H�v��0�e~��T�ޓ��%�e���fYc'��N�֜�B[�PJ��������nQa���h�� N��=ދZ�{�옅o�X~�~V��{�,�`%�(��&����V-���&�r
��@�}r*^#N�-��D�Q�1� �(cj�;�)*A.�v�:��Ly.Rg�{����B�տ�L�����Yr!��E�� ���M��f��)��[1���f�2�-k}��q+�'�]��29���*S��[�陀DϜ���<eq4�Z~���{���S-�<i|��Dc��u����H��Ȧ[�Z�'#8�\]74�d?h^��޽'�����P!\����3arre�e�>�Sm?q��p�ė���Ǭ��9��Ӧ�*�KN�3¬/L�%A��HEܳf]���m��'ӌTJ���}��7Nݪ�֋���Q0kd�S
=Lx5/�碐|���Y�6̶�y��?�4�P>f�,Ѐu.-�"�f\�?:�q�ވ���A�ܣ5Ն��%?L�.�N�����P$���~+��t�Q7Ex�d5�d}�#�C-D(Ts1�Dڦ�1*������H�J���s�?k=,4l�|P�����9`�:{I#�����@e�[���)N4�w�^z����Uf5E^��:�W�7�tN� N
k}_��3�E;S�V������7�<l�`,�i[�� #:�D�,��yi��'��+
�>\?��K�8��&�"#\B�O�3��2R,^U�+ci������I�h	V�B����Ex��k��s���K�/��V����6x\�	��[lFn2먶���'�n!0�]�ᓭ���u�J>�6�q�L�j�8� ꍻ�D�
�4�c�BȤ� Z�m�&ׯC��򱰝�h����Q|�S�V��3�ODc���Pfme��M�ܗ�6'
M�B! K�/W��y�A�%X��)�۱��;�i���O /t��JF�Q��dܗ�XV�;�[CY!u��O�P����ʹ�#��ቧ��Z2p.����$�L�|h?s�CTy�ӗY����>���g�vX/�#�O	\�Bk>ϷZ��r���6��a���#�7��Q7c�.vK��8����}f��^7?Ǔ��,(�l?}ƥ����t�t9I���������sU�K�^��xv%��^����qc��u���1�.s��?��wh�<!D��̖"=�Z�&EX�H3�ѐ{j��Kz�t<M�wrYp�ɝK��(�5üM�ܶޱ���ºB��Q�q�j�u�l@���/��,$�؛I8>?�y�9f��F��Dr]�_H�9.��V���gMbOJ+���(S��y�A����DM*&,�7S�-[����X���0�Y�c�ފQ��jb�ʕ�"���Ce��d��[�s�z�:{��n<otm�C�wɡ�T|٫��Չ7�+1J�����^�l�[�K2\
�v�Y���^��W�$X��E��,�}9��JϪB;C��|�4k�:�)���� ��{e'��S}5�{JjKLm�e����%Ȟ����g�f�E4q��}Գ�"�J@�������)���3�	�b�;�c����zvm���n�os�H���{����Z�I���̡��+".����fR�\@���R�t��ꄣp*�Yu�s���A�A���}��4���V^�z����{8����"�_G'�{��n�0Y�����~m[ @� J �����)�pͧ��O�WvQ����!�1|Q�񺹭g��8�cD�-_m��f��)�U��*l�/b��م�X��iY�DH��;M�E�]y�SI���ŭP��<҉v�g)c)�ʫ*v7Q\S�`��?o�;u]Ī�-��@n�KS�Xg~�lr��x�*D$sO��?�,?�`��V�`�Y�B�4;M����.�����,[�����Q�y����:�ay�*��.9;
c���E��V�o�ҭvG)�uk��	uu�S�%����=H�g^�T�+��%п𿬓�߲8gĪ��TnFv!w]���Gҏ�r1�L�C��������,�v�S�s�����<�H�b�H��0\^�j��!�fk˫cd���;~f�0��TC��<o�4�B>�P��1(8��ב���{h8z�ږ�����9�
���-�s��G�u�,�]������Y\gϑJ2M���ACC$�����9׻>e��V�8�&O�
�.1�%�����a~h��|ѧ��@R�.�[H�A�x��cn'`)�HJ=ޱ�[%���t��Fwn�e�=����J� �lrf"�b���'~�+�d�_|�����*�L@)�L#ee��b�������m��K*Ie�5��خ��u%�Y�ʽ�z�?�*JI��5qT��iq� oۅ�TJ�b�-bE\wd�g,����p��$H�xV��cb��ٵ�$n�FV� ~����Ob��PňӰ�ǬH�d�Q���0� ��ɋ���m1+�'��A���Qù��h�d\n�L$��Vگ�2�֭ Cۘ~t�3ܫ�T1xi:M*ń�$Jie�>/�����X��80�
`�Ѻ�&{G���̺���{��Ā��g){M땂�"��̵�[V^��#�U��^뫙��׍G�Q?7�b���@�Q&��=�~��Ֆ`�����\�_�����\z0�j	�kV��V8�hw�_=C?�%�:b�$��>�A���""�tZÓ�����(S����fXN_N�����*��º�Yt�6��&�`Y�IMt�-|2e���Qӻ��Q�N9M"
�RU3��&�N�����'���,���aL��ֱ���wp�7,�r�nd�WOv�q�-�eu������_�ے�3��{��T�����Q}4Nkㄻ��6�y��:t��f$m�y�d�2N��
����-ശ5��CJ*��9��_�>+�����hlM}rF}p�?*J�h��ʇ'`&���)'�q������8��"Y���r�8�~`�c�|��r��|urW�G�$�A�計<��{EK;�_>�k���#��N��f���a���:���ƫ?�K����;�-,�;��� ^��;%Fv2څh����r��<�i�=�8���+e�X��h���t{�+(Hr���t���E�sm\o��:���$��CB� �Z�@"Qn_��UU����,�QE4F�`8j����M�4Q݆eS���ˊӢ���\kY��҄�IU�J\06�j�W��C�Q4^k�آdmv���f5��PA�w̗O�{�A�'}$�Se��`Z�P�97T�y�\͂>��!<�VX��Y�·4c�XX+���+��� c9���ׇ;s "���'��b���ّ�:t
}�Bˊ�[WW�C�M���T��q�r�Đ{�L�p�`P�SXw�h�rO�R�
�޴X�,7�Ѱ�8���E�..V�͎��p��w�]���y�o'Z	U�
!��
#Ƽ�lM�Q/ܖ����@u��$ޤ�}�)�tc� ��w�+S��L�����s�\��7��Rh1s�n��CO4�u�X{�|��c�8�U5K���r�ݸ�|�nUH{qt��W�*�_�K������)��������ݰ�L1éCC�a\�$7VX���k{�I�TI�dG8.�J�����AL;#Ձ��$:���&�.��\��m��r���/⌢�)y?L슕�X�&���2��P��3ehR<DL�#��췍'k���0{�9\�qE�/�`�~ e�)?P.�gS�w�&90Sw�ۖ>�83�R���� 3��?��a�n,���af�"���
�����~�&�2Ƴo������LR���IKՏ�Rp�@|s}��OSNJZ�.�*3�9��,t�-��P#���5�n/���.
#��@>u���t�"�?}[����ؤ�H/X�Lh�,="ֲzaz�-��zn< w�kC�Ҡ�[)LD�|�m�,��U`-#:�퉩�@zx��T)8�U@G�%�Pqa�R�
+�� �USTn�_r�,�4��X`�7E���/�Nɖ��Ԯ�����&��2$p{:P��h�I��ܱ�3���}e���g�n�ڔ�}�d�5�]������Yn{��@]$/'�36�>��(�P�L��׏g���DG7�{��ϑ	�(�Akm!fmyj��5�H;~����e+�I>Ej�ܑ�Q�|�-���<y�gĖ�؝⅓��/����\9�$��2���M�T�v�wK�N��r�:N�E#��(�E��5v��� ���0�Q
���Z* ��D��7����"�7��7̓5�@��B�#WdZ���'F��|��<��|��ayc�v�r���ޫ.D3Q�i}�6�D��XlxVHYEB      e7      a07���Ib�ێ�#i���!ZF��u�����^�t׹c%�h^D��N_���~Ҩl����X����?���b�����ZM,3�h�>�`�-� ���;��Ͳ�T0[��|2��lZ���Ji���N���n.����u��>nk҉y�5���