XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ml>zƐ��c��T.�p��D�:p���І����.�]�w�9��/���j�E���c�T����m���u3��*�:�d_MPv��%'bt�]'{Yn�f���
	0vj��[ʽ��9�6y�yr~F��8��[�j�p|:m�.�_�b��/ �r��y\qvE�i��'a^\�'�sWۃ+��fa������K��T	� _�VLW���i�\����<�Q���p?�B��7F*>�H�-ƫ�ڎ��Fd�����{��w^b	�Rv���r�cd�����Q^B��šq}��k��Nǭ�P8�z߸oֺȠ�W��\�� �j�Q/��nW.���f\ܡ���(T1Ú�����P���~�2Fr��j�5j�3��^:}��AҢ:ΐ�w6����c��D։�-�4Eǿ0��R��
NXc}��V�#G��Jm��<���b����"=8�?�ɐ��T����pC�<����6�E���@4g.�݅lm��6�
�W41@��Ÿ�
���&P0��@6?iD�4�_T!�}�N!���^�Kq�N�>h�nn:��g��V���m+i�(?���o��z�[G2&�d���P�e�Z����BM���K��P�{�ju�1�> =6����랿_e�+�
#a�^�U�1�kJ��)�c؊��`��Ʋl� ��b	��n��\ىb������C�]1OP3}�Kq���|�ӳ���������4�+��g� `^��I�u��%XlxVHYEB    c763    2600R��g�(�nƎ�F�es.�+�r�X��C�K�	=�/�z5��=͒{���p�㭇ɪ�2���ٙ|l����Z����KR�nä��E"R�_5�n�W�����V�-��-w����$A�x��\n>��s�����<ح��S�0H:d�_6�p�g����TԐ�<��T��X��~����v6�i?^!���ImI�#�/��z�d���m�G AT�5'�8B�nM���u?I|mR?[	00��rh�#R����#��a�x'ia �H�VAjFVd.`~���s�-!������URuĽ��٠�?���[Y'}&�S�|+}5Yl����J���<�2@+|AAQ��ZSB5���EKA����Q
*%";@��Wʨ��Icp�2Q7s�����_h���h�ч`�,χ������]L�/3c���Õ���/BH�h�:9k��� ��>��&E�6^O�J�� �Q�9���v�����'?�9�y����?W�(f-R҉�P�iήZ�(X3��%�+ڦW6Ȓ�#%DڈrK�
p�P�)�2�c��om`��>u��xR��~������ӳ>��E�o���/뙈�ژ����D�j��,�[.%VS�
6l.��dS�'K�(��S40�E�w^3S9ǩLe_>P�u����p���Z�zX���~{)Գ�x�u~�l:��L�TAI9IV���ߔ
�VھlJ�&u���~������!;���4�ۍ���}ӳ������r�G/��Գ�'���W�NT�U*
)��d�L'�x3�刘���`����}Y�����y��8A��4_�b�lҎ^�\��@B�M>[.r�a�l��������q���e��!�*��}\��g��.���z-8O
�r�No�b"��-�V�˛K�H�������(R>��t����#<�m��'�h[4F(=j>���x���P�!(X��z�`(�� ��E�|��A��U��_�h���_������'?CI�L(��	ۜ5u�F��΄nq�D���%��B���D5D�Ა��9��lN2����L�@xiy���}9�|ZH�����=�>��U-�m#U��{�]���A�1۲��G����@E��+.4�s�j!d�DD菸Fia, Ӿ�'M��eo��f�m�����'.�G��L�O 8S�ܯ��xM�a�(8�
	��)�CH���a�OQ���ꮛؾ��33�͚!��)�"�۴U�oY�@XS�  zc�F�.���;O��Ԭ����;�l'n5|�D����t��2������� ��؞p4����a�]u���W�����p#�1Ő �5��f˘�F�-Á��,�D����6Hā;X���"=��ށ���.e[Q1�i�u%�������i�4���we�1�ԓ7O�<���Ǣ�����y2a��P_�co��n���%�V5�����!wgs�}B�K�DҚ[^t-�[쥕8YԼ`���30A7(�e5�*�=��Sy���/ʽ�j�q�/1�x~(}��\��dZ��"�~.tU��~+�j����D�<�t�b�/��<��
�m��˝y��I���H��O�ExoydU�ݸQ,^v��d�.pX��%v��mD9�5O�0��4y3��m�6�=x�1���a��ЭO�kA��2Ka����>P肸g��[)��Q�	t�V��oD�_�P������K��b\�Þ�>-��h��g(���!~�r��b�sg�?þ���\i�ˎ5�ͱ`�pyN���3�+� ���]B>ऀsM������^8��Tv5�j�Ý oT�N��Vr��%0��4)hD.���^g�S�\�즑+�K�ro9�ĞN#��l7C�@$��F� E�́������P�v�(�,�-��6��zBMT��S$�ɴ�ZF��9s��oS8�r�7.:��,C��:0(1nR`�&���ˠX̢�޶�t>�4%���&Lj���B2N��z�޲���I��R�yC��&�cQD�-eږ�^�O��g�}���7�y��
��{�^�RTb�K��j���i��o�,�~UQ��?��/
U���U�
v��ZY �">����^�tR8rW'�O!�'�F��h�[�������ȍ���|�m�~�"�߱�e��0j�ە�����rQ�	�H@zbu�8&Z"�E�K�;Ͼ�h&��լJ��v��Ԗ �L��z�a��eט ��AW)O�!�L���A��jDPϏ��
	K�Nf��	&n-Pn}��k��X�Ȱ�咲��������P^����$�_-��'m;7��<�n�Z�Y�C���ܭ��^��k�։�B�n��١o���9G��(f�w3vo�m�����s�PJ� ��%�2������y9���W�Ή�6-�<AW�^�#�1��ե,2��&�dsd_�L��#�>�[䆈����vo�dt��Z�"�ĸJ$�/���į��+b��3'm�n������6/~�w�tƥ�[=�52����Y���/�<�O�d\�M���urp�Bu�tlc}���˩$,�K�[�^^�߫�Y��=�G�����!΄��׻S�-e�vC(':�<�A����ۖ�sb�r�������7z���e*`
W�<>tШ/H;��D���Μ+��9�[��-�Y�u���Z�~�ǁm�V战@]h��{��)!�fK��o��S��+)��	O3ٲF��υ6J��j�(��؁rnc�<(x= n���u.q�4��+��}���,��	�
!6o���8��;��E�94DS��8b��*�ZB��CM�������.�C~���/kY�T�(�f���p����$Qe&D���En,��~�ܧh�s��V+��������2<2��΍���[aм�ࠍ%bsw��w����s��>X֓���_C��(����/�e]�w�@��V�]`C���"xN!ͼ�[� ?G�<+��W��L�X۝+騙�k'��7�����9]a!w�o�r��!�D8O=�����#
v=@�O1�0�7�L�KF�ي�E�E� 9N� �VTA
��J"M�ݎ7��v����f0�K���a*X��R{��l0�FZ|2���5K��(X�	h"��.���ޯ�Bd{(&D��c�+�����|*�8*���eL6?˛�$Ly��X�Z����E= ��7�q���G.W�����(	�A� _�EMqb^�X1(͈�ǒ�HC5��JP��q�݅g�*�����x�(�����6RK3��z�v=�U�8OwR�.4)�d^��tc��p����}Qk����������Ӎ7��T\0[���V�֪���/G5��V�Of�c
��5b�nĵ�IWE���_`<�b��t��z�ʛ�n"�Q3�2�uVXE��i�"B�`�u�����QJ&��fo�Q�shn"����p��E�~j�����1 t���'
�єD�bɼ���ќ6�c���'��'�y��x ߼��xsw��@(�P����j2���K��7n�i��yn��8�&C:-%y�RK��'��A3*��f�?��w�_�o�U�����|i3=O;�
�P�Y�>p���2ж�wz��l�z(�<)��~>!�C������EƩ�	�� �d��I�&�v.d���Ҕ�>M�9.Ʋ��sV�El�hQ�:�f��uw��o��e˿�v��b:�3nNV���ӽ[QI�0�+�	E�W�ХQd����3D�&��8�Z9|�$�Yv��!PJ=�G���K�[;�pzb�\Z��K����^h�����i��='��q5�1ڂ���~��Nr��ם����[r�������{�$���_$����Gt�-�� \�$v]T�dm�
��5�H���bؕ��k����k�җ`���ltԊ��|��C洠����{�t+���X�JV�v��~�e����=�3@�]A�\��:�����`94��X}���ƺ4'�%<b�}Ŭ^&����
U���D�
=h�!)�NY+=��i*���*��C���:NeI��!��A1�T �������ra1��dU@�G����m.��J����_R�u=�oX�_�|jС(������AP��!P�d�a;�q��A4���5�ă=PR� ��,�l���%w�Ir���D�N���$�Ju4Ux��(�3GV�i/�FyM
�C�rqy.&qY8QU�Ϣ��i��~���x�v��H!�� ��Q���\bM���J*_N\ਯ�{1Z�`�.�-E��W{�έ����f�����s�Gd �S[�ޞ�]����a�>a��/�x%P�Pr�j����޾E3U����ss����2=��A$��;��E��]�r��QWw�LHm27&������2zo�"=R[�o�.��e�T�we~���C��5I4��x��v����h��jWd=<�� T���nm���e㧿r·�L�m�����l0x����%�@����~�U��Z�qGf��d��8�ї5�Fa*�ǻWa��1�]����T/����Q�X��� ~c���bS�Lj��:�׏d��iƐ�e�t^f�Ǫ僌|���ךF�3�|��$�[��T�0F�s��-�?sZ6�#�=�#�{��/Sg��W/����s%�F�����Y��߳ �GQB��_ܼ���?��h��b��
��?��f��Mp<�v`ւ��E��`	�$�y�S�i����_�=5����$dt	<�k�c<��g
s#YB���k��|�S����:��3�B����o�W�D�Jl�8���/�tIZk��xtQI���%�$�>[N�u�S4<����)$���������D�o{�����Y��c����ρq�����Ř�ש�+W���Nү�_�]\�%
���e=ض�lb�A{P>�N�p��:qMaԎ��뺁1'	���إ�m�v�[�d j�jW:_�O%�������@pf��ԢfB�!_*�'CMB�4(<�EDBGH}�LJ���2r,���D���r����7�����/����D�þl�wFXQ�J��s����y��X�`�=H��6�`��$�iND���j9Η����A7㐳��Qt��ybi!�@��4�Ԕfj�BX�0j�Ǜ(<f�~P;��
S�U΀	J�_h�=~&L*W !x�r�2�-�
%�\��T�)R�����K�n `����w;-��L�Kwy��<*i���!��sV��pa��Py�6��ZSo�]�R�L�!S�w����˰yD�,�!5���
mr��wb�<I�D�!`�x\�nu	�T�����(��k�`�a�J�bޞ
�̪�|�]�|�G���М��ʮt��J�k�k7�̠��(1�4m�A����z<��}��L[��bnC�4��DB?�M���xJs�����Z0�6�gz �?�|P�ޏٯx���*�l�֧=��}@
���VP��=+���UX���Ӷ�'>�9���>����@W��ǁR�lΊ¢�G}�!bx��d�����9 ��Q��`U��N����6�S�]vV�G��b�}4�!a�)0`�@ԧ|��H'D��ё�����������o����>@^��_���j����q�4���[/� c10���E�(Ub�����_u>�|I��.�M
���d�&]G�k����r}��r���z[�W�i�1�?7J�ǐ��A?�� ���/��9hRg���]��f�eb�����	g�=g��|p��Pz����,qlF��(*�{u�}쬏�Q�,����8����C�hkA(ƽ��T�:\q��ub$�����
+E��.$���[#���T��*�TGE�E	"����B୎����c�����������P(&]Ȇ����X1�
ؾ2R�'��%��yh�=�_u���s~�x3�~���f:��z�۽H�f�|�����av'���^D��=�x5�X�_A�M�m���2��ɰdg955�!�	�͕"���$���a-1	�ch%V1��A'q�^lG(*"6i�6��$o���,�|3/����Z�-;}�L���?�̓��G�ۄwN-D|Р��X�l�6�3�F��5� ��i ,�K�*8�!7g��~
�O�O�eW%��>� �T��Ζ���\��;q�R� DV%
��*0sEMUv80q ��j"hM����8�'p�X��N+P��b���^����S�=rY3�=�g��;�4�K�C����N����88�����W�Z�;�>ud�?�D����$�#=`T%�G\�6���N�mc�R��Y�.k���r�ɲwx{`�x4���qr�T=7E�;DY"f[��òT/�LV��=�uv��7s�+�9�W�e���M�/X>��#{v�[d�I��j!�P(R�~\vN���X��<q\�����yS�7I48���Ӽ����HB��M�3C�q�d�k��m�I]e�a�W�K�<}6��Z�9�d�*0s�I��ZՅ}��7�_W�V�9�!m�"q�Iئ���uI���:�?��Kh}��>t�R��;P�=2:!�Y��6�_"�pCj�fJ9�[|?6�h�mB��M��gq���%ȣ�=\���v ���}X^�A��4�X��������6�$��݆�?hy/&���P�}�Q�ù�-;EG��E�_O�.�u%_TP��~i2�N���܁���o�5[��U��7xS�Z���9�-$0LJ)�D���?'�ML�l��2W����C�j�l�A�]~q�l��],�C�`�gq{c)���[ v�k�m_'��U� ��T��e<�4YR���i��qmۯj�&��ɤN�Ȃl�M��Y嘥������0#���!�q��ނF�Fl��2��MY�v[
.șxt��aK�>�&��� ?�����	gc����nΰ�d��zE �_�ѕ��+%}���R�iï	}��-�R����ܹX��*8�>j��ɜWE��]�B��Ӗ�R�LNcf�όxj`�W m|�S@(�U��m/������N��"�C^X�ؕ��o2�7�)��'��N�D��������o�A��L��T�s�CH�6E!�e��9m��{����s��W���jM�F�2�5ӘI�}�%���<���e�T���Q��bp�3[��u�7d%�͘����=�"s<�������iQ���b?Ky��fb.�vE|�ߺ\�!K�ֽ��g�M����Ͼ��c����O.ߺ��i��q�mDI�ҟ<�������-,4��8Ή��Pl����F�q��RyV��9��4~2h����%6�<����2�zF܎1� 0�`.~�;�c��� �B�fC��
#�R��u�J��ں��ޅ��^�Y�XJ��T��h���礿�5&3\7�֘^�g��}��pG��u$p�F��I!uA�]Y����5� �Dx�,��W�a���\a��LG�{ݻ �%/*/�vƨi^y÷�z�e�|~�g��C@| �Ei�nA X������{�d�J��ӆ~sA��V�U�=�Rl�/e��w�4>en��p,��1��O=���)Y���lv� ��C�&�<��U��e��|���r+KkK�J�U�sA�ear��Xmwzi�'�rxe��ZaBkC(,��抎��n��ʍoŉ[ĉ���hٚ4��I�#{�%��Kp�- �#!��]�p�@��}����˪��6�dl0Ә���^+5~~����$�t�_�a5�vk�!*m#䭽+��͌�|o�����*�>��I���]|�?��;�1��8��Cߘ|5�{292��G2��D�2�K��{��غ��uN�A�ܹ�g e�������	.�f�������<P+i�]��}!ͯ!��IE1�/���j�t;���c��%�f;�U)�^ߔ��}�����>�����8F�NB&K�eó�~fEv�+")�<c���a��5��7a�\[F��3�j�tҗx��2��S4aQ���[r�ձ4a�hz��	6�Z�l�ʩ�߆��x�>h�a�1�Au�g"���E�,�����ն�>l��0���VF%�����4n@%VkkA���y�/�z�"���-Q�>,6I潿ײ�?1�sW�4����\ӿ�5�����1X��ֱCdb]&BP,�y�zz�L�ᡀ��-�פ
�,	��<fZSkE��v��� :��Zr����CB��.X�Ac����.˧Ud�JeAx� T��BlQ|\m�1�hV�|��%J����� �8p��`�<���v����n>�D2��;<���b!��Z�Ŗ� �+���09����Ѭx]��}�Z���֠u6��\'Hoσ�O$Da�[��v�\�:�fmu�;t2�����F�|����r]��B	i.��%��Ҭ��C��j��X��B�����~R�Ѥ��C�ㅪU}�l�|�NI0I��1�Z����6\t ���-�s�Q�ޝ�+�b]���g۫�$����{�>� Ƙ�,j�=��t4�JxO��ah��:K�z�Ė�I����gy���K�A�8~���(�hz �-�*�t�ۀT�|��y�)��������nf�/��Ev��Q)���ܑ�
���˭���nś�:<h�^�BQ�E��/ƺ<����g˧�G�3x#ym�hS���ưp�����I��Y��^Ϛ���f4׭q)��]�ѧ��9�b�ot�q��f	]�}; ��I`���4x���M��< u�q�@f��v��r��z���l����<[i*g�F�m�P�9L��K����<�i����� ����`Sq[��ʹ�8��r\s�o�5r�4��s� kllgLn�I8��b�T��1�)���x���xf��,o��K����V����>I���jVD7�N�_f(P�V�{-��?�ѕ�` �UW
Á(K��c��Ei�@.�;@8�r5> tc�s�Q��5a6.^��vO��k��Ǡ"�+�@K���S�JZ/ƪҢs3ޱ�>,Ƥ ��]d
1���;��d��ѿ���D<U��d���KZ��Z�ga�"��� �r�䯆U��_d����VK�-V��0+�Ԫ'	��M�M(?��k�;e{R��{J��`�.xߴ��$Zy}��uRw�J�:���}c��)��݇"#���c���FD=��(��7_�V�t	�t�֭�?��àL[�ɁF̸�����8!�"���`C�)� ��F���`�!:17���	�A� AU�oM>-7�yt��t�-�:�չ<�N�l��]��x|��/�N��Me���s��D�$�=)R>��l3Kz��a*D(��d��[~�S���'��D̀��fU*o�^ٸ�i	�yx ��¯Vi�d��\\h�H��*UGƝ/ ]�2�+��M��y5Y6Ϫ���Stz*�?|�u�h{��m׽0��e섆K�`K��R1s緺_����G��﷪��F�"��5��Q��v Ғ"}��vW�2q]d�8aޔ3�M�Z�#3
��Z���
g	��*��_wf�8��J$B�g`