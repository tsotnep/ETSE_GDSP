XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iOD�:�������\��1��7��<'O�z��X�h<D�ѫ��	b4o|T�����aF�2"�w�w�w�S�̾�zf،�&�C�� ���Y��B��λ�F���
=c����o#L�3̜3����8q���o%�y\#������8ML$�}�4���\�3�67�Za�~;%�V�kyV�?
Λ2�I�%��b�}�m����BȜMඈ&A�o� �J���Ǝ���h�`�F�.QYM���q��L!���r��cU�tg�F]�=َ�p��GA�d���S���ցt���-F>�Q�Ӏ.�Z����n����*�Y<��<��X�,�Ͼ��=�����u�mʏb`EV0Z-	m����bS]���O�%Β$���2���a.����$)���c�Xnz���C�r$2h��
�������D��lLQft�*Һ�N��V�Gy%�#�����R�����i�뎶�n��!�#���v���`�e
�lT.��Z:_�8�뷫6���%��R��Y4H�ԙx�6Wh�	����=���OC׫�Q�� ��ݍ�e��p\�D_��/���K�!Y�@MD��WC��m?SJA���Wn�,ǠD�8ӼEw���&�\��R��:DU����@%�T��$C�wF���?�z�C�M�<Z���P%�e�w�*x:�d�^���35C/'v���I�!�z��p��gO~W`#��\Z����E��]4U P�����VQ����e�LDܛ��dGdB٥���XlxVHYEB    ea93    1880\g��P�R��Q2r�P�yB B&�ۮ�g�;�%@�~�fe<:Qc�Bb���&3�7�4X���	�A�-pu������0^��W���6j۞W�#W�!��z}p/��^j|���L�W;��.6P/�}�-��l�l�`t�Ij%{����=:�p�F$\�v���q����3�����ᠨU5Ɔ�T�ۢ���绷4(��0X�'��@+V<�r�/H.� ��{�������T�q����@�D����oc)
D����S���������M�.Bԉ3!��K@������:��Z���V��]\�e�8ZXG9ߟ���o$ҭmg���m���f�}I�y6���6(����	`\�i6��U^�)�k-��@�ݥ&������ܿ*�o:����,��h�Y�
ƅ����lY��T1��U����+���G�}^!�^F��q�'�V#4�Z^�����꩒z$ck��T���2�{B�P����M����!�ťB�y��y���C�֦-OM33+���!?T�����ք��Q�����O���P�4�Db��e��i>�f�x�6�`uE��}�qL_�l�_X;OYSO���`��L�Y��S�\��t�%�Xp����	@Е����w:�f<�:�q�M�~��h(-^v��%�R
$��#��Ԧ�� �š��w�t��[��	�eT���|��`��'�6�Hɤ�*�yl8���G�{��2+��!�&0����Bø-}�l�m�	�!�V�a��.�~����Z]���������ɫ7d�N�V���۲*:��nYSM���Q��"�ЛY�
�xk��fX�(�S�cs,�����v;c�N �zF	3^�='�J6����HF�+��AAQ��d�����7�P���-��� '�>�h�2EIw
�ۇ۾�j�;Q���i�98��"ڍ�$�naOz-��=/�:��\b���8�)��8��I'���Y�	[M�a�<[��ڔCn��i��2�����<�H�SE��|���$��p�����S�c�!��
�W�9�O썎��D�q�c�������w��'p�&�g>E�:Y�]o�U�����֚=������c9Op6�yHQ��"U{�1)�h��@]�;7�6h�,fv94�\����3�/s@85��Ƞ0Ы�@Z7��L?�I@��G?뮬�_���M���TW!z�x�83�!ʧ$�e]e��wKh��f�࿔����R�Y��V���E>��p�w/�I����.B��^��qS�����RwJ��UNs���������dW@��"?��<z�Pw�?����X��'YR�L�ﮀW2��,�y�Ι\4��æ\��(��G'�6�9�y$L�7]��Q���46N�\UmC�U�Q��	�)��&I�^��S�I�
�g=g��N���d�� UE��;���ޛF{���<�"����u�3�`B@�ĺ�D�)���[ +3I�B��^�� ���e�-�%f/���q��\g-�҉��5�`�Q�a|{�Bx$+8���/��F���P[=t��As�9?��|u6[<�_�5�,�A���\s2r&u� G}6�`;�1��Fʓ9����1��yQ0!�R _H���A�qՄ#�i�A)T���[�d:��Is}!,�)%���_�E:�o.̹��=��-gb��lKSǤռ����p�9�M5���V"0O����k����C'��>WusO�=�K�e�NQ�Ckk�};��.`�5;吀RH0�j���(�mǨӟ��Ø�|�Zc�֥�Q�r:�#L���rx*�JGA�f��0xD���C�̹�̗�'da�礆픕���fF%�`�hY�C�<΃yɰ&�/�e���>DuTpjhq��OL=�*)_�:�e���q��~��	O1�.m;zQ.l��������I.)攄kf�I��[���N����ʾ�U��}c�]��.��5gFk~��^�X�e�S�la��;�651�I����1V5�
	�0Nlwg 5'AL��C�$/����S���0b��9�Ǩ���^gbI7�IK��2�z���Mf������ L���IV�%����G�a��	��C��^�z���p�W�ę�s`��\��E�^�1��{�nC ʴQDcq�X~��D���xv=��ŷɥ�b���H�u�V}��B�6��#Z���V�0O~ �Z���fv�y���r!�3���wS�*��G�u];[��\Gp4E%�Q�N9���u���L'��:�U5
�P����x����*1���|�����������5�q$ഏ�0Nk����k�s �7����2(��ڸ�^�V��#fhm|�#��ge�E#�P^*��x����Eh��w���Fك�Wh��(��-��:|�l���7=����92\'���C������N�M�u��`�Tn[c��1Vy�3[��]6";�� uj.��1rS�"}��?6'�[��Xq% ��@�ٷ����B�@�C1 ^��bTc�d���X�K�_:B�'V\�h
�����/8!\Ӡ�'�-���Zp���o�P�����1�*K�����p��@�Β���2��?q~[#�������[�zaU~O�I����ˬ�)���a�u��8��w=�t
2o�Ä�k ��7s�w_4>�!K@���A���	��:v�K��$><�ut��xj�6�=�����x�D�X�kv"�<��8�$?�e�,,�UfB�����VYR��Z��������Jۑ���zWF|�p�� ��s�Fb����ze0!W=q�˝�wF��t�&�ĪRu�&�-���^~�M?��da��۾C!K�/|��,�e�{�y���WV��]�V�ڕ��>��j��x/Щu�u���,;�f��v}D�z��|Ƶ�������6�zΤ�O�eB��C ����h�`L&�����V�	�5�f7��b�/u�VP�7��R/�8�/�oY�:��ؼ�v 7`�ҷ3���	%=jܵs� R�[��b��2ڲXgQ��j�*%�__�iM5e�g~��o�+K�^	��:#�Bi�zW�&~��=j��^V(E���
����z�~��U|e��	Gq�QV[KHOٓ�������>��Cݻ���$���Er!p�İ��	�mؼ60���l7bF��{�U�޳\9���8k�a6�2�'�b��j�BfdМ�B�(t0m�s��Y�bW\h���3���RP�����p�P+�L�v��~��π�;�f�־�Q��]� �?�}�"������ǣa �@Y5�4
"�(�4(I����m�q��h]CG�Ǎi�z4�� �b*�*�68j��b��<# ]�/s#	�n{O) ��7��Μ�p��+lٲ�瑱�X=���A��1�V�=���U�8@{���-,�,��&����c ���)X�ue�i����1��B"���Q�E4{."����B>��?��'�KfU�:���:�������l�1�|,���~��Y_����Zhgz	% 
���&����<����ӧ/��Op���=����P��I&)��z)�{��zM��Q��A?�c*'9_�i��Kt'WGM�Rb
��?v��cP���RҔ��#��	.��
+=�>�͎,�����Jf�!l�i!n��)��'4��6M��,Jn�
7�%�րy��r�)��We���tǸ��Th�E�Ɍ�:�85�Lfg�'
���t�JbEÁG�u��'N۲NnZ��u���N��[b'*yL�bX�f�ވ;K9�XA_ �>��Ttz.��㴨�Yu���<�q��iEո�/���5�Qc�9�i�������^��ɶ�;�=���Ph#�x]�+�E�G���K�����R������]pԕ�s����Azs����.�7u,�������ډ`7��fD��h{"kSL�$2�g�\�� t���/0p�B����yQ�F�Z�ɺ��Pٞ��<��2�{'v��gM�㭻�+Zk��ֽU;#��Z��o!�t;��B<7eM��p�l�oI�Μ��::��r�����0swT��B��`� �'lt�xv����R�o�U)����,P�w��нI�����0f��d�e&T�&j=��-�M|����.Ľ�,
�7�����6V�� 5T�G ��$}D�~�4��5���=;�$�p'X�k��$L?��At��Y�Ҫa8�}$�~��o�����������!g�3գ�4g>�1VR�A��&*��i�@�"�:5?+��*�X�
��w �\2�
)�PpX���M���(�I�!� V}��sW�C�.qd$���-J��	4}�4��<�Ev��A�=����x.#ͪlc˻�� E� ��K�� 6�?�ͤ�-�ه�y�( �p{2�'���Ұ�'�1���&��ӎ�d;I`�~��0��m�Wd{ҥ9����\���^l,���;�7ּ�|��Tg,:T)��K�q@�l��>(,<������4�;�g'�2�2®��vX�e��ț��<�bz"N�A{b������V��g3C2� ���U���˅ժȼ����~��G��YU�m �1��է
!Zm%>r:�Չ6�r\5G��{��e�DE� �ߵX1�0�jIH4x�e~ۯԎI�ʮ�Շ�,g��y�\M=��?c��'���B�{'|��N�/�L(�'���0�M�ذ�:��m�GYx�t�Z��L���8�$�b'5�R����߸B{Z��3�i�dm��!�M������Z�e.�H�:Ō�����Gp_a���Ѷ�e�B�W�)'�Jf3��i������U���%��­��~[�_����k���H|y[�y�E��N�����\p��2��u��#�<S��#K����'P�=�Qu5��� õ���Ajr�W���{�\	:�<o�g��QGX5�f�R[o����t#���S%މ�snb��-��✭�j����5�J~pC����_vN��#�P�T�3B�?��P>�2��)u��ߒt&6_w�Gn�0^�r�0�$C7�e�=lO	��}�k:��G�,�l Ӭ*��Ǫ4����g��8,!'j9ɜ0	���� �E�yFJ#po���L��^�&�,p [����1���.�sOa��S5����p"�eRA��C<�-B#�.���<H���AO6�/���JF�]B�`�E���毅Q��U�ˡe�B��f�Qm���d�ѯ��"�=�L�'c�
���[K��*�z�Д�%����ҩd���e�<b�5*��(>�f ��9�}.Y��ff206�#v�p�����cTe2�q`��":��x6�7��\H&g�����~�ӈ
"A''>�$�Ol9�������'�Jcz,@.��`Q��%5�,�G@h�a�?������A(F��u�e�.�q�M�k������X� #��Lw^I
 2!�a�����u=�W܋�K�	�£$	ٙ$Sa���)2�{�%4���8dIÔ��4�"r���VL+l���߀D�T�ц<3�^�&��c�F�π-���5<0?:�ځ\%�V���䵽JP�ׅ�wL���,u[rRJ
��)���>/����'U� }���������s�zQ/ee<����V�f<@�j��\ ��O���#�Ż�l���U�#��e�39M�K)e~s$r�d_��R����b��Z��Eһ�aJ�!ʸ�CLPz[M�XMN��xC���D���UR��{�Ek@s"��B8A�E]LN0�zq���f��L�<8�h�/ɼ��E��r^����(�ny���1)�3�37��A��~�� y�QDZl��84R�9Q6P�'�[4 w!n:��xG-���ľ�M[��M���@,��vGێ�^p^�ђ~�O5������x,Gcu�ڦS��._��+�.b�9�z�X��5�K)��l[Q��3h.�Pa��	i�HM��yT.w�1��ՙ�{�KF=��7��,u:�5|Λ���j{�t�՜�pHg���ā�XvHu]��$gd<��o=d���Ԣ%�s�A�����O���k�����/#�ul��Q�T�WC�ϴɚ��i�-����hm�=ֿ�q	ӷ�z�