XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���h��:T����J�����Z��+R��7߶���(���b����$�O�E!(F1�N�w�z�9�;�	�:�����VzR����G����oW����iO�}�� Ԭ���c2G��w��\�je<o���p���i�4�+VAggs!'�<*��m��8ARGs�K�ZK7���B9��;���C4;�
Vl؏oX����9�F��Da�H��F͇�X!|��^����K0OWk�A���q>��b:_��ڐ�5Q�KQ߸��T|��1X� O����9FĔh�L�y����0P?��ux~BNP���"D�Լ,��x���8�!W�Zf&� ��A���3M`f��6P�ۑ�_S�{b:fh�<�g�i�h����2�GR�/�����*�a�TM@�ByC���f7',���1��䌬>K�����eק����@?JC���Gu��D��6'p�?m�m��c{�o7�YQ�;<�A��-HV��&��c�CyF��������&�����d���Ww	2@���{Sߟ&R��S?��HmN��V��%�u�]�>#j�L2MĐ�7a|��)W�S �\��B��@d����n��f~%r'avX�&v���r��퀭|�Uk�����X5�ڠ�dse���w�L�F���Ѣ�퀭ʆ֋H�_N�"o�N�B;�h�=�F_p�ZH>�N���=��P��u1,�qo(���q���W�hR /ևg��4����X�m:}=��Kź!�b�p;\9XlxVHYEB    162c     850�e�,�g�����J��gŦpӟ���L4�ǧ�/\p&��,ʌ�g������*�<��L̆#.l�8d�ٸ� z��wˍ/%��g�UJKۼg�NHI������eS@&Ɗ��F2҇�`�8.��:��P��N��k�B\c�3Kے2��GZ�q�	�vn��<b��X��D�|<v�$/��B�Ƈnu�Yl|�c|C��oi�l�.Jb��W�2;����H��TӃYG�!dD�3_�xl��ǧ
��Q�l���z*���t����=͘����M�K'$��E�� E��+q��ӕ-}HR�wm�	`E��0�g��4�Y�l3W\�[�|�Ťf�v�u���q�w;�������	8��W�\�0�9u�n�$F�a/՞Yj�=�n���#��YJ0�]_/E�Y"�w&�b�1u�Wc�*��E$8�f���5�-�P�2S�N��ؐ���R+g���٨�5F��=h�_-���jɥ���h�2��IT����� K�m!����P�ŎX�@�'��Q�>|�<��ؐm{x���\k6�2v\�9iZ��Z�����D�}C������kr�\���|���f�]�؍��[����O�Fc`��i{�*Y�i%��M�=�T�r
/��k���l��ǻT��`�?�,��{J��5��X�3N�Jf_a]E�x&�^��Ԧ�6��Eq1�����w�hX� 譪�+5̾�h����2U*E�'�����p�����i&<����T�rpB��N����
]lV��	+t�2\��D�;�I;�M;�y�0;Vo@��@Wҧδ��[{m�,W*��5肟�<�p*��8%���x[��yc�hM��&N��'i`���O��qu5��?�u��v�T��'-�cy!�	p�r����
g�]滰�lX��rx&�ń�M�| ���E�:�	��Qc�B��[��蕍�T�� ��mC��(�(:O�a���t�#"���淎��t"�v�IˑF������emk�F���$��{�Ǹ�1��G����O��H%O���¡�����	�q?#Ɔ��ч�1�K���������ad*t��������wV}�;W���x��<�c�r池Ŷ���^�{��	<�K������b-na����~�wP���x��Xk� }<����Ԝ��a(*H�uS	�P<u��מV%-���jn�8NGQ	�N���0�0;�rD@t��x^�~�u깔�1i<��1uV��˜w�8GHH��6��u6�ur�S�"��P�{M⥘�S�|��~"�Cr(}�0]2[H)����P��d�%���s+���||��>��T��s%
���B2J� �c Yv���y{A��Z�`�@3���E�x��o���oµ���'v�f|�`����# ˦jUME�yؒ5;��ʭ��
t��S�
���_�w-lb8Ig/Qf��L\���	 )�<jT���cJ&�A�����v�N�?��)	���őG瑭�V,\ K���;Hr��:E�O��s�e�ìݲ�s��P�y�R���H�� 6�����#CV� �ݵ�a��ݍz�G���C�/LCY{�5K�.Q��ͳv힓U�;-�kL;�J#�tOŸ�ͩ����R�T�׃�+�,��v+�{"3Aq&�T�W���Z�&��ʵ"�D�I��?xV^�U�=�e7ۛ�Cű�h%գ_J��H�#\v���qی�P��̚a�g�̺XӉ�,W��"�<^�YP�q�<�!Kٵ��Ӟ���D¶w��X��9Vh���}y/�	o�1s�z�����(@U�s�e��awaA�����Ά)������O^L0�}��_��<|Jh�M��-n�[�ͣ��j0���aS��W^ڿO�\�LG#ή5��`Am���QI��A�K�8^�⛗n������Ȥ	64���E�R4����rX�\�sO�����R\!T=<�P`	8�0��y�x���>�l��r ����^9^��ӆ�4�%t�㗑����|�@��)k�~��=W�5��u���ʭ�Z�хz��ʙV%��N�G@98ͼ2��L��c^���]W,��;����W��(ȸ�