XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�L�ѻ!a�Ph�~��.��0�T �O�&����8'qn�x���#�K��J�g�A?�����A�Uᜱ��ƂoX�K���ǖ��0���#4z(�k#؎��t���C�{�Ѐ=:@Z�i�<���n9K-2�[Iᴘ����w�KQo0�������&P3��ޏ�ᓙ���R�W����|q�˯Np�������z�y`�+f9-�aD�n=0$�E�H	��O3��c�S���Q�Z0��ז]��;?Y��l�ʤYѯj�4���bf@'L;����~����ӕl?=�B�֏q��e��@y�,S(�3�-�!�n��!���vL��
S���Gqe^~'�X�%�T�Z.[��Oc�����̜G�g$}�\٪ٽ��2O���m�0�,ߩ�����GqB�I+��v;oa����qH��*��[�J�����Y��ޔ+�s	*�e����:�����	)����6G&bJ�N�,��������������t�G_�d��W�<| s^��lEM��A��8c��'f��V@�߄�R��e5�vy��J����#h��Tʾ�k�>��� ��4{$��gg�e]I7�;um4���\��P�������Z&P?����{B�=��+�7qo;�/R&rF�� `�s� ����<�c^�:V�`}F����V��|�=��ߜ����"3>!�G��|K��к9+E����9�A�H����;x O�j�2$Fj��&�%j�t�������/*�b����ۙ�U�Fʜ�XlxVHYEB    fa00    1ca09�Cf��C��k;*+������t_�9��v��;��B��5vV�bH�T�N��1 6�[��a��+���0�c�X��޷��M\h���h}z2i	'~��RU�������e�7�@�C�8v����5ծ��0D���z+a�����o�݊8b�������B���G�XV��l:L�w��̃�Q�],p��ʐ�GW?Vo�x��`&�8+������/��F��5�P��:��5fG����)����Cy�b�qZ�W<ZըgY|ۢᑟ��&R��c�7-%?v�^����,L�a�$V�p��[���X��y���[��.G�	*��-�fD�i_f���E3��è+�Ⱝf�Ǥp��5{�mϢ���F9ΰhk��Z��*L~\����y�ll>�8�^��fEڄ��?`�{�%��ߒ|����mw�]��ȉ�X��n�"�a�1�3*��jFǺ�+��ϐ��� W����w���1�5S��[�ʗ�E$O���x� �w5�ŀ+8+j�>�sZH�Q�]�O�I����XE���'�l�Q��c+�����Q�����k�<��D3sN�2" �NB�f@�e9���^HT��Hj�nW��8{��z���
��n��{q�ll--�::x��C��������������l��q�SXpg��J]�T�)14]������.}�^����Ǭ��I������T����K�gB/ĊD�aqwي>jh���R��a��Ny��*��u���X���}lO����l��3����¡*q�A����ɿ�"E�b�����]E��Y��8@��;H@�M��ޟ�w%�7��,S�`�"�FMt���J�ܡ��4ׁ�i<��mF�t<
GVa��r�M����ǵ˘��4o�4�Ŗ(��?XƐ�KC󡽷��Zđ4�P�^��\fӂZ���cW�Q(��Kn��k�I�'��Y7bvn���y�@s��
i� O��q�m�o~z����z�fg0�c}�O~�!�����9�e�Oo.x8>8Rf�I � 8v)���������P�|=�ԉvU׻OL�i*/4�(�U�3eC ��Y��|��e��c鼍i�`fͯ�VՏVR��D�A��`�9
�?�8��B��N��o��q�Fsx踆�Ve��4�'ڰbaӄ}����$l��Ӫ �����L�� �����Tإ,�_b��~Ǖ*䍋��*D��z���(���dI�o]�
�(�/��ҝ�r:�}��z�ʰ~�&�/A��C������r�_���֋�3��IS�L�-t>�uv�P�C�#��L���?�ѱ��&)k��Pu��.�`S�s��%~56:����'z+@� _���{�K%(7���=���2Q�t}3�L<�}Hp�}��	g�?t�����Q��	ӈ�0�����R���[�׉�GU}+���T�x�2�n��/�B3L�C}.r����`OGX�e�m�G�^�c��̻_�YҼ:�ef�V�y��-���`� �h��5`:��V�!!cf� ������;���z��U��ykL�D:~ʨ�D_�ݒǳ����VӰ4tz�_��^�*'!$�^pG���_^�u�)OA�FȂϿvM����Ү�c= ��K���y�y�ty�h��$x(�q�~�d���Dy�ZyQż����:��죟1Â��+��V�Yx=G��Jo$GМr)�;q��K���
b�^�.˽W]i�.\[2�oz@�5�$� z�6cX߂,�E���l�Z���c�j�U��&(��06
��B�Xp7k��*�*>a�/t�jr�/��_���]>1��P��m�������ɐ<&�%��=�F뽁��dq�}C����\��5!CM�>iyR]���w�j������P�������߂���V��r?�MHJ-T��xۗ����6��fR���]~5v�����:�l��>�+w�b�p���z�g��c���8{Z�����֠�d(��_��g��2>���7s^-�����fT� �ۢ#C�`(��Y{��ʿR���^�K( ���_�=,WM�\�s ������ ч��
�wˉ�\�+��!��R��W&N�A��� �䧞�*C�o�:�bR�����O�Rra�!���]Zmy~���F?�t��H��pz=�H�O�r1ϠZ�����Y�k}ρ%�F�"B!ϋK�q��ٷ�ߡm_+L�+�Ev��7-��|Vd�s�M|f�CM#��y���8R���q���bSj`?ל1���CJФ�K��/Q��ײ8���c��$��-���S�Ԗ��G����
i�J�$ꕓ�Aڍ��+"�o�#un�P���'@4so��%��R�'�P��ϙu!��"����������'�`����G}s��R��?@P� �[=������a�r��S "��=�%=�a}p]��ˁ!Mh�.�	
���jͤ�'�Q<Y����Ӽ3��$-�F8�5��$GR���jD�� "�&>}u=X����b���#�I���ۀ�-�~s ���zL������÷�T�I�,$u���Xd�����p�7D�mQ[�c���D�:���K�Y���]b�y�p+F��*�N ���Q�.-�8=���n�`P���v/(��͗TM�2��3���)�%BZ/��(��!�T��+����'��\��ȟ�@��n댽�=W����y2���AWYq`�E��k��[��Nu��:��-K�N��>�Z_`�5o�AMm*���&O��p�ܟ���� ���0��y`[ew|3�J��vH���q��-O"x(��|��u��!|�ݭ�U���ۃL:T$7���`K-��+�a��� ~���hĚ옵���r����P�qpꄤ�aځ���h�d]�C*��'l��gެĖ���+�v�aB8s�!F�mģ���8ֵ#B�&pRZ]%x�5I� ����/@M#���j^�D:���v��
R9���CE�w�0�c�����K�:�
p��Z�W�;׃���p��P��|C�')�y��gI��\U��^��Ik5{�ql���q*�z��n�;���������fA����l.I|�<�8|��1N�׶�\��E���H�#tR�^cx�;��]��L�S�c�xYvi'V=�eC�JE�_�Z��w����#o�|��[P��)��Q���&2��7ʅ	ؠ��!�PI�db�� �0�O�lw�'L*7�W��;��y������j��9�����g�L�ݽQd7n˪a���l�~e�o������f���S�-�@ԖvlGg�#?� r��-G���^��I�I|�l:C!���{)�j����d:ӈ��=Ƥ��>��k�qI�2%��(�sa�M�ɋL��.Ĳ�D������k��
�T��[K�T�O��:w��������Ăf�����O�)�V�I%k-khBH�Z��-�]�Ԃ@�S�F@b�,Pȴ����i�#n���{���6+���`GCB�,��y3�]i�p��
�;~?!O^^��j�Ro$�'�x�NE�ٽW�Ӧ�i�{'�(���=�AJ]�����l��Y��O�(+� aW���s}�{�V�.+�9��ݱ�o�E�eќ�(���I��g����t���@�1�=Hh2�!�D�ߥ)7V.*Y�E���d�=�1)�Nͺ�4�#�r~4�C�En�-�L=���?��]�2�<�rTsF'H�-O�F�����}��k+�߲k�0�\��v���_x�qP��C�g|�{�q¶?~^ӻ�@����9&얊X��Rv��~
���3je�K@$$Q��7��8��ax�B5�MuT','Cq�i�s=�[���#��T9�n�P�C�2���
�;T��R��w�AL��Ͷπl����XR�H|U���^��C��!�.�ވ-��03z�HJ^7(�qoc���՝�ޚ9�:p� M��$xIFB�Zx��gn@��xK���e�Ѣ��F>�α�!!ϊ��d�� �A��D(�`)�{��MUXN�U�_	r0��'3���6{2��'�l�]8z���IWA(�Ǆwq����Ď�-?j~0pdE�5�z�0E�F�kx輽.{ڠ̀�W���[���X�:����rU �=����fD�Μe̐�-�oȨ.�8�����~�=n���ه����i���or88��7�G��J�>Nԗ^�Z��Txs���#y�9�:5.;��oʫE�dd	��=)�`���j��+l����_���Yxf����6hU@��vE�������ܤm��g�Kx#���^ң�Z���f��S��F0���5���7����59�R�i�n���cB���K�b&x�
��(�G6@ߩHv����v0:�m䡐��C�u�W���/��cu�!�c,	���=yt�n@�@�W� �]��r�{kG(�|V����z��9�;��ib�AY�w���>0�*�-��Nϡ|XX��K[`�����ٲ�����[-%��R6�MyEܗ]�J<��t5�#�}Y(��O1�l���+��lD2B]�ŃD�<�/SD��R�seV�u��M�H���]g�I��I<��>vn;�R�ϸ��4����YX�d��5'Xj`��K�Tp�>T)��ƁR���?��q~(U�K��ނd�/�+�b���pk�wY��
l"�B�):�*��K�"�� ��[ \`9 w��p���eF�1���ؾ$�XA��ˍ/A1��W��� �3<A�q�E�U_�U�0u#�bG�h��:�%L�Wd?�8*��w�v#�V)�=���ƤajHC�ɵ֑�CA����l���']��)"!�DE���/	�IUJ$ʑQ�g��*E�~����x���o{�b`X�
��Q:�?�^j�q(j����>�'�W��3#Z�)�����Q
���k�ѧ��b��o�/��0!XQ=��T�Q#h4b�1Ve�u
"ξt�? 3h�)��R��u>�uY/�g���*}#�:��E�!����E�J~�H���*0"�l)���Uȭ�!	y�f�pՏ���҈�S K��-�Ktm���ͧ9�L����W���s9^hO�Y�ӳ衤�aɝ/�SP�!5��OuV�{d�@*�M��>փ�d7��8���6���x�#�Ɯ�ԮB���]�$0��@ΐ}t��m!���^�K�E �M� ���c�W��ә<F��Bh�}�L��V�*[�?�n�I+��x9,_0ȑAy���q�+4�3l��9a��e5z[QlY����d���l���r�IOǗİ1���q>�*��;T��8l���V��Y��F��ͬ&xց�/8����c��y^ZE+�N��%ȋ6D/T�?����� 7S5����L2��������DӅ)I8��f
���Z+*,����C�r�N�P�Tm�����b.�7����b;�F��z��*���ؗ$�A(j�M�]��e���}*5�t�OE(�s��\�x���WHF2�������������r���R�>��D��*^Q��D������*y�ѻ�~�4���
�|ʑ��L+��3�����&(!�s������?�S=T�N�1TВԸq�n@;a??^\z��;�U�CŨ�z���S[���G��M�ja�[�;���Eԍ����\>�O-�j_U6�����j)w 8;�"�Zǫ}G��F�t7�V�
E��!r���j%�Kߚd��BxM�hhI]��H(A>@c��G��k�paPҗG(:�t0R�{V,U
*@I���{�_%�̕��c�e��DFB;N��@����
���q��]�}�|W���x3��z�_�$��gh`�[��N�><��cn��;kq�<���l��	v>�g�sO S�P�@^o(.jodW)�JZN�)�M���w�cOi�u<<䘬�!P��V���_ �s�r��nÐ���!_���"5�.�":�n�����p�lm�*d�TI![So-t��j��z���Miب�u�9 ���L^�8���3ns��C�<n�~�<�W���l�1�
�p9!��x@�&�J�y���� �F�As7��i0kvXn���@,� �쪋�HL�}jI�=Ǌw:�	\y��nKkV,���u����0��%�>�z��C�dep�$H<�%�8�F�~��a$:���=�U���D���ԫ��`g+�k?u����2�8pCQK*��.��:�f��Y9j��|U����`���K�h�-b��B�1�:����]{��frG,!�!��Kq���6Xp,E\�Zm���<���Y�Z�0�zf~��;�ՓNYy�F��܂��ߓ⏊{�����8��L���De�e\�?���4[�)��:�A�m�I�bW�Gk� �p[�-2]'e�)m�n|�Q�N�9�l��=�Vİ���Lǔ#�ّ��	S�dbt�JyE�u����M��N�N���PH���d �u���-��`�g�Z�C)_nb���{�t��^��"^՗ח�
����U���(����y;D��Yb�g#�0C	o�Flu�M�O6�A�Gõ��+���]�:�<���8|iS�h��D�s�G8uS�ay7P���;�i�X�����b�j��<O1�9���u�3"����l���鋳z�Z��sj����o�|M�K��.�������.u��F�~�9|Ya���/�,v�rJ$v������pﱻ9/��x��u����g`~���S����_�����4�Y|"&���e����6eD�C8!�q�Z�|�	���2}�� ��&H6ԞG*(�zo|�iq����M>4��{G�CK�<2��ٛ���S��}�,0��j~�[��*�d(�{��OaGٙb��G���A�8Q�~ŧ��*��2�Y{0��^_����0,����\^I��~yʐ�ހ�&(?�0��q2��W<�b�u+�~�;����*��@���p-����u�sЪ,���g=DJZ~颎���t����|��~���pQC���u��ٚ�.)�K�k����D��7*��X�f+o@�%���Oqj�L ���pI8�7D4��g�5��Q�1�=Z�N������Ϧ���y@�ID�@�1��\j�#�~��mt8)M=h�(27�M��*$�Bр<ڠ��e�pݡ�Z���N@�nZXL!c��q�B��*�מ��
��9<.��\��I�i��?�s��R��\CGO���zsOʉ�d��?�?0�F�Τ=���Ȼ�x�b�:ِ
a3{c�b��l4cWS�C��B�=,�XlxVHYEB    fa00     cf0zo!N���z��꓌���Z�a���a����~Iy.[�%+=K�*�	tP��8� ��uғ�K��e:"
�A�NT�[#&j�mL������X���Z�	XھyW�u���c�j�9�蟰�_:b�;�Z�t�Z3(>��Uh�F�発���xe8$GE�jd���ͧ'L�I��#ȅ�%��k*r���{�`��v*�84�$
lɆR��Qy���NIg���v�w��mY3�i?����̊�Q@-ӯ�eJ�v+��9�N�#ȼ�R=�L���b�u���A�<I�q��W����^X��k��Y�h���R�$���显n�o؄Gy	ե�(����@�g� W��S�2�R8XC�ѭnwh%�-\��;M�_'Jhi�3�	E�)*���t�9�y1�u����v�S���9g�j�ԵΛ��dP�!�F6c욿'��#��O涿G�<=7�7&���ˬ��p���:5}���dW�%�������!�ut�{گj9�*'��W'J_�!���b ��j5��ȄҐ.�
y�p�Q��9���Ht��*��tA��Y$>�t�z�f*��D챽���)�-�=3 ���gW̓����G�f�[�O�u�]��C�q6k��J�!�BU�o��	��-$��?�3M+M�G��1�7R���  �R����w�q��R��<<l�c���C����L���kB;/����F�]��{��tuʽ�|[x4�g8d��R0Y��UNo_���5I���Q����9 [!Kd�ޒj��Ba���FJ���S��fы�>�#X��h�a��C� ڣ,K���<`�QF�Z��e�g�����Go�2���|$x��d{����~բT.��p��F+'gn^�imNi�cݠ�<�QqJ#�L&��0�V�o��0���
���Z�vc����}����K'�u�I��v�K*A�U��_O.�e˓hʘORѺ�pmH�l�ԋ���Z��;U)AO�|wA����m��WyiNO�`��{��1機&T�U���\�{����[��}Pȱ��z\>�f�0��Bat6�v����j���M��N�P�N��q�?����Ԍ�Lܣ��m���AЪ�4Y�]�p#���˔c�ȧ��7�Iul�������b������fE�MY���:�T{Ub+5f�鈶��*r��%�ge}��M��r���{�ј����x���O�b�w�s0�f45���[���dA��͸NH���e-�e|�32d�����M�$��r]ʅl�\9W��*�0��V�g�.-���H��t�`�ל}��D��lW0I<�|U��ۤIQ
bo��@��	���6L�2lU�v��#*��t�
m�=�ZM��sR�vky�f
���1U�5������|�.b	ZFD�� �J2Nv���H����%z^wN��t�򷥞�'���Й���"�^~�t Vm1C��;���m�R=j �GM��_#M�T�:�|@�(6@T�1>�wd����P k��j�ȗ�^�P�hi��I`܏@����N�y ��4"��'J���w�ٝ�.�J27�֗���_~�u���?iQ=�?��e�/h*��v8����l<��A%�ח��hӳ�jJ0�"}��'%���,#�+B��ݲ����\�h��m*�ܶ��p���@H}�ͩ���ت�Za�jH{�� ��+�� �}5,;$�!���,���de	Z2|t�ѯ>���/�����x�>��j?z�r�Ǡ��l��g
�]Y�$��Ea~pJ9�u=�ez�l�H9�)jLId�Z��=�÷���@%�Z>��A����F�2
����bG�s��B*�p�m%ĖբTG�~O�rx�z��Em�D�8<Eoc&��������YbO���y�-�Z�|#��]}�Ve��f�ؐ˖�T���Rז*��a�(H�[ ��8V(|!3?sԌپ�s&u̼O�yU��j'n�~������^����@�?
�mG^&�P_��dH��f� LeyDs�>�1�m���h�*\���:(3p�Z:.����}�f���<qT�J̲���o�Tē���RNC�?ȵ�C��X�ݑ?��^C�!w�����Q��IH����b`ڙ��]H�@�Xf�b�'��Q�_��E�*�Z� �l@���j�b� �*�`Տ��I��6k�,U�^խy���b���Cs#~=��d� a7mǐC_�T��f$�I��4�e<К��_1M.v���`��! ���L�o����ΰT�|9��l�,f/�!�T�N�G�B}@ޗ-\{ʐ�x�տ�^��[ؑ=���[�lļfK�[��� ��i���nh��*�uj�`�ћj�8+��2���P��bv�^�G�{ނi)?����S�)t=��5�v�v���֟�����O�x}G�(�5W-X[+<;,@����]}n[>m�G�L'���"�y2�O=�������Ӫbm����S)��N��\�	@�g�h���g���e9����"�e׋c'� �]|G9�D�OD̷�k��~d���f��.��_��o �g�{w�d̏T�E��/�)�|N�|�L�������TYO�jQ�ed�4�Z*���g��_DV�	��K!��0�LмK�L�2�عj�pUOC��_<�߬���$jάX��TUQ{�{D��u�i9{�E�	�Y�G�tl�{�̨8�H�1���.���1*mr.��aA�6(L:�ǣH��P��C�N /t�G(w�~9��1����5ˈ�-4-A�����E�=4$'�������fh�ӃjM� ]��x2��Zw�3��i�D���Q��}
ֻ����j{�o@ ͖�.Ko$�3��J��'<��~��=�q������3-�~&;

`)�V����
��߷#|�	�E�L�/��h�����}n�Mݳ�6��5�a�la��._�ڲ
$ZR�KB�((���%nl�!g@�,���)ƪ�� ٗ�R�j �iZ�&Eo����p�NI�mO��������S�K��u3-�Y�M-zc�&���-OPf	].�Xfn�w�����Q������O'�Ji�O��y���1�d�yS�".�|~߶��7/�u��<�����T��_yȣC9�y�{�דpS̬.��djVa���2oz?�B�=����U.���6r#�^�^�>��{3]N�K~�X�����g�4t��8���0tF�\=��E6��J��m)~��
�Y��\nXlxVHYEB    3981     4d03OO�5�ouo��VY��I�װ�$�hU��`څ��A���_|,3��ce'�L�F��޲`��V~}���!�� v�KRv��zr~$W����'��d�H�y��!�pM��r�D�
�Ml�v��쬳M�����)f����ڰ��QQN�X!�'0ضKd�v�q�4Nkأ7����/���n����w�226��b�;�Vd�S�qB<lD��Y��ۊR��b��USH��Ui�ίI'MӪp���K��������y~�ⶀCG'�4���%
-{�����fID��{���9i�ׂ�@����� !�q�5Rq.�&|��~���V��V�n��#u�tc�����e�a[���k�r�~����%D�ъfb�)�C9��mw���	fw	T���:�L���<�L�Wj_ԋ=�c�G��Ԛ�F�3�T��Fͅ�(���YW�|������N�Íj`�zt[lC��a�9���!��H��ܥ�����E=5Hn�0�SH��������Av��.�z�u��}��D)�Y�D�d)*w�. �U!���K�fX��xߤ0*���e����+ٕ��;2!�bfLkl����������ު��@5��9�F��T�wA�N?I��cډP �����~�TG�CQ��e$��n����]R�����%�b�Kdc��lsN���u��J�H���o��"�e�m��v7��nk�OI����84�@;ZJ����5�tŠ���������yR�j���n�p�ObKe�4�r�Q��m4).��@�/P���u�u�kE�S���.�����̐�5�$�wO�C�b���⭢��.�<)<��!�i���;p?�L`�w.!w���
�
�l�#��̓�k3R�O�V�/�*����ݼ� ��YQ�զƄ�d<ST����8&Ua�/��3/�m��4��y�8�	[z��4�h½~$�P���ݞ���!�k�lhԬg�q�7�$��������c�ib.�������Z"��+�0�}w�u�#g�$�ˢ�����>�������lkݛ�;�yfv���;+:zL�G�u��]�KPגWqc�@a^�A_fjLX1��Pȣ�LfT�mЗ�b�)j0�6��@��B��XͰ���u��h_����
��܀�4��U�����Z�!��N��p�XB8r6�8����&^�Oo�%���