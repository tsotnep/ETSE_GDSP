XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*y-�	.�,8!�ZZ�[���*4��}�ޖһӞ���B�Jȥ�a�$�Z�r1��LBY�j�n�Mr�-�t��}?�����f7Í�?j����"+p�YY8�ȼ.�`Cx?�J�=�xP����	�e������	�l���R8}���8��џ۴{鴮�0�{� ܷ�j��j^�@'<�d��g��K��= 6F.��.$z,c"�3��E��*���|�懃�ȥ@��Nn3���_���^��7V�C	L�l�ݵhX���6�5�_FiS�V�u�w ��0I���s�@�ߣ$�i��Փ�z)�N�c�.�5�L�M�'�Zu����בj�N"�w]�'~�q.�`o霿�CX���<TW����*�"�P
���oG]8��nB'5�|\�'�[b^���%��ҽ���
�9�V~�4 ��;���Ie�b)fw�8������SN�a�X�d2�"�6�A#�튇R\.���(�4������V6�u� ��9��J!�щK�3�T�S±�Q�z�F�+�r�<�����T�~�΄դ� ;�W���(	��>�;���@v�D�4�_��o��6�7�Ei\�������ޞ��@�B�8>BNΉ��^I���]�gN��@=�s
��I�䛄K��z��+Dl%ճ������$�bĐO�C�[��aG�"G�4�3�"�H�Ǵ����}�>J�D�J��~��z.�f�s�o�F���88��;1�(���7%'��[[S O�CF��'"�I��ǖkXlxVHYEB    3042     c80f�Hj	/:e�0����5ߎ\VH�N�n�;ų�e��j�b���'�5���4R:c�.���Kb�zS�I��-7[�>�@?�U�R�9��#y���8v��z���R�'X�j{Z���{�|���!o6�3J�J�����jR����!����],�����"%�����:�&�o ���B��r�+]��.;o1����D��M������Hvu�,�t�۳���y��87��^ ����,�|O	�o ��㰜�
���	۲pY2�Yґ���Z�EM�e�����w�ׇ+��M~�V��ƍ�L���Wm!2�(�r"�|n2H�II`��rj�����џN�/E`�,�V�'��^��S(��Z_!ɍV?��[D�w,i������c� E�)G
Β�����-�h��{�NtX�9?c8��5ci/��(: ʧ���F<X���<i��1��.��jE�Q�E���6	#����V!���<�g�u��-!����:Z-���c:t�̘¾4� }ˑj/�D����g@�tId�F'�F�cV
�O4*=����h�a x=J�67�D�ddw�<�k|��=���&�����ς�:�*��k�u� ~��N#%ߊ�0��T�޴}9>��l��ћ塖��]c�Hչ�1�ks
�60�_qC= �э����TXj�jg���zy�;λ<H�z���Z0��ĢN�K�!��*]��{#���ۍ���+q��k*x`"�������d���jF$�i��Y�6��e��Ŋ#��P�#tvi�7S:g;�qͿ"���6����r	E���I�R��ĭ��[}e�o7��<
�*�W-��ȑ�;���7�,�C��u+���Z����(��k��3��/N�S.X��Z7c�L�]
rvf&�Ou,���-9K(�!�<`J7��s�$o@	�5��w��dk�͉袨����[�����8�|R�A�wd7��0�x��çJV	9���i�˟��ӿَ\6� ��bN�޹�m���<�jO�c-��A}�N�?��2�>=ũ������R���[g��q�"Ͼ�[?�j-���?�@I*L�������㨙BHz臭�]�sS�pA7ePf�-�[W\��coB�x��U�L��*L2��Zi��0L/�@	}���f@)�[�+#Zѣ�_���"�8��vc&�pbRJ��$�{SƏ�m%Ul�Uy~�XL�P�׽�Pԥ��,5�2�܂g�۴���G�P�d������

�[6m/��g�^�ʏ.X�f�?!�F��d3��*[�]ԈA��l�����g\����̮��8�YK������^�r�*��x:�N �e�)�����"h˖B�-˲q�^�P�ގMm�NY�lF�N\�d�Y�ר°�Г�m�x6���ry�'c����7��j�󰓥�#��=�"a�;I���e7I��0t�4R�($�ʄ~�d�P�� ������Z��������6�L0����"���l]��=t�UF��Q �QF�#��`���i�����"��*4��}���H��*h{�R�|u�BL_���5n�r ��tf��2�'f.ڎ,��;�Ɍ���5�0]���pY~���)��,�y��d�Z��b�
8��6`:6���#�@��4�J��ʹK=ܮ��@"z>�&��X��.���aP��wKSv>&$�ϔ�h��
�<
�8k�������x�k�ڙ#�;Q6.0�e��-P�WL��gx|VN��L�0�*q��WC r��d�9Cϝ�Vuޙ���ܭ�-��;�-d��0�X�u_�].�Mڶ�����k�cՋ�B͆&���q�`���)-a�`dޢ���N���?�	]�?w�h<���14�*��mS,W�l&�=1��^/EQ���Ty�hMd�`���1l=#��t)?�ȇx�J����AD\��@Qhc��.J���(f�C��Q�������#��ƿX����+<�0�S�ت�����q�&�I�F��y��J�}���FiPН��ҙ��E�]�P@��x8�n�����Zmְ���WžWv��v��2��*�g=�@1�L}Y�C���-l��=Id�	��q[��L���Aa�$�@���ɽ!S��Q��j��'2%�׬�#�ր��L�&ݡbs�c�>��J3�7gy���x��C:P���ȍ��[v�>W��Q���Q"؝В�����Uܹ�����J��KO�з��$�Pi���w��py֝&��FodB9\�d�KZFSO:*֝+�ں�ӓ��Wv%�".�!��M���:��M��7HYP*���ֿ8߿_/p�zf�~�Ş��J��W03���Q�������i�>8��@�>�y~�]=v��v��~�z��
��Q꿥���e�
axeuc��(���0{�	ʹA<l���M0���F�@_3ZBm���0^f����Y�0Z��������I6$�����,C��.=Z���d��S�yK+��J$��h'df+�=	o3��nW�KA1&}MNK��Ӡ'� ,����sð��K6����Q�gDT�h�Y��6M�0WK��0� ���!K�����}�g*T�2ƫ�`�!��� $2H9y�眹'w��FO�a!���-x��J���Aކ	����do�����[o��¼5T�c���	��	�u� %���uC��@"9��Et���*��� |@�ee%k�b��ăI�e�To�c��8�4<��d��] �������9�
��ƶ_���*Np�@(�k��4�L���1�nȺ}�a����|D�	�/�O��O�ZY{2%2���qRe|�S!I,1�gfx�}��Z��icRM�i���#f��j�	#��鿌C�g*�N�~����`��;� oh��Y��3LST|�_<�N1*�(�O.>���l��*5���b�PS��m�j�f_%5����W��/Ő�-�ő��,�Տ�%Z����e6SjeUw�5�b�5/��[XL �o� �J$���.H����;PH�將p>�u�<?i���֓8�<D�T��S�)���H���3iu�e�i�^�v���9��ʱ�%2�X�0�F0�������no)C��d��