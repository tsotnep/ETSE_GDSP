XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ip��$$��F�j�����>��Sj�Ph�dua��1�Յ���c�">do�,��A����,�n�q���-Xx�%�f˯�_��+z�Dr&��i��E0)<�+�{K�Ao!��/���}��s4�rW�L��6Ӫ,;��͸��k��_\d�D�qF�:������35:v�7C�=�w��Ω���>��ՙ׌,6��0����&�t�VY��]�P/ֻ��`�D�}Ya`jIz����X�$�&#�����A��W�2�=R�xhŇIs��
�����������0���q� ���̂�����r�1��;|,5�:O��!'o��ה�F�=ۿ�41�NX��ɜ��O�q�� �=%;���' �p�rر.��xJ�pPl������,D��J��F�Z������u"W���k�o�C�l��Ur�N<x����k��(�GAC�`
�����`W�����ա��>ǵ��׵uӡt��ǵɹ���Oϸ����Ha�U� �,��-�@ۓ�?���ε9�[�ܓ�b>AȡyI�U�t��8���{T%A�266�	�wq�a����~�Y(T��Fi�V	{Cr��	)�4��:�R���5��)��6P��r�������A�td�피X�0Q��zh�<cȄ�_mE/DY���������ڭ�`g�6�\ґ?A�4�CB�U��d�-�^��4;Q���M����*t�z�܂����e��Eи��������o�z��q+R�#�7�gu�Fk�����XlxVHYEB    b631    1a00<�r7l�R��n	��U(:�3�/
v��v�9~�~�B���-����gк��F�G��a'$��>w�����3BQK|��p�j���C���"����±L-]L	fJ� |^�b,'\$,`ʐ�A��_�n��KmO`���$'5�����P'G�Ì�i���%����n�h.u�Fߞ�6�x|�$��� ꠼&�xc�U�=����NTV EHf+��b|�0c)
�>uk6~W���O
x���n�d"�_�!���&!�"����:���Z�%~.�\d�D+�����*$�[��)���Ѹ���˞�s�9���.�P呈a��E\
�|)0X>��A�om*���|�A8����q�J�A
��lm�p��B�����
l]�g��7��\EWN��W�-���u�I�3S�Pw�d*�E(�Z^{��s ����v�,d�2�,=�˪w��f�Pq!����T����uU8�'�|L1������\�[8ۧ�'s�p���2<��s�~f�O˫s��;G'd.*�0fyW�>���#�(�p���Ea�`��41��b�
�?\��#C|DG�S�t��}�}���[�7����ȭx^l���n|>�"��t����b����MbИwd��E�������/� U�f�He��˘`����e�}�h�E����N�Ԧ��uŨSHFE�>�;�J��	�7<ªws#V̿ ���p�-1%����[��̔T��N�=L5��y��,��]U�-��Y�����0ߒ6�i���!��uF7�GBC�-ld�P��#�7±�cuE��5?&@ⶔᐧ42�����Yؿ>��𑘨�BGҷ*��?�5�m����ƙ/�G��m�~��y0�*q�B����¯�x�F�s�۫�p�I�G18]F��I$���ٕY��'�������Y��m����J ��%a�
Њ����*u��k�.���z������sk:$t��,���l�C+q��a� ��V����f�Ck��WJ1��t�j<��8񓻞����d�̓�1|�a�_�g����Xٰ��e2sf#�&P@fou�,c7GG�cf�Z� ch����#�
ͫ�X�G��}����F'�W�1g?w�se�����hp��cm��`$�S�ԕ���`�րo�
�L�Lߑ1��Ȫ�ۗd�s5i��\�۸X7lv���B���
��)�߃E�6�K��Lq8����7��(�c������;.��3�ф�����'QG.�^Oz�d����o��FQ�
�i	-�V��pB>뾴��G�Us�x�����7�v��v��M��Ι�瘘`*d���K�e�����VDc�I �\�PgsF�e%��e|�6��J��1is�g�f�X�������f&�Pz��A"���&M��Z�"M�yiX���X&g`��,<�?�]^ٟ:���?��5u���SV�7:�
�����^0F�Km�k�~�2��o�Tn���N���/H9�>T�#i�D�Gc�׈L�lA��旧�BeAG��p�RN�vf8�F��k��O��-�11�*�O�-E>�TU�
�9R�ۍ�k���A�on�]y8�Θ8���C�02��KD۱�O��{@4��O�y)�V��w<d��?p�n_��V^�qy�[(5��k K�|O~�&4�2�3oȎBZ���>N�:Qn��ڭ��_7�L)M��X�q����Lr�X�G�^������
-�������Џ#$  SISkŧB�Ȩ�Ϣ�������^��B�Z]8�:�웥t�G1�Osc�v��۸@X����˴[������G("$n,~'�z�A3�]�
�;<|����y]c��*���C��I^2��U���l��z:�� ""��&�U4�7�}�	PJ�Sf��^�ׅ��(@87/�5����v�8���޶���?Wҋ�p~| q� ݣX�\�Q����wE�,pz�y�����H��k��^*�S��iZ� �Ao�P��Ɵ����	% ��[DS;UQI�X�\��`� +x	8�����v?z&������x�J�����VX��W�*�O��o��q�iy)�ʉ�	ge�dv��ed�������B��`@9�Q�ھ�(mXSPK�`/֣� �%�F J'��Ġ�D���|�#���eq�Yw�ϩ��
n��]����Ho�L;yy���
�F��J�7D���O0O��y�Gr��4A��r�;]U�"sG�:9V4E�Qh����C�Dײ0��֏x�������K4�b�i,��Zn��>�u�'��@?׽�� � z衉�N%�n��-a���ɍ��]�*v��i�Ň�͡aJE����vv�{��C`k����v��� ��rﯳ����z)�ܨ�
�T:�3Q�����Z���X��9b�x�Q��VZ�
�N|���'F ��N���gkGP��Z�
ԥ��y��/��7�7���F�T��t�o��H}�L=��&�~D]��Q���
���ޔ*�����w�1��MCs�\�B�#(�`"x3<+a4}c��ܲ�$Ѯ��\�C�H|F:`�����r���L@�N�^Rv;M��#QĬ#2᥆{�P0�[[������;����
�2�w��x7A�4B̯�W[�]a`���@��_C�i�f����d\�;m�Ϛ��<�Z+� �b}D8�����!ƨm������|���)�[���a=�����"�-?EA):)�_ƙ�{�������`{1�A���#�F�n�������ǣm	#W������j����|
���F��F�@��I��W�Wf���!W���N�^�ˊ���r��p׺�������l;"5�ޗUCԭ���Hc陟a���{���:�.V��{��������>�Q`��Z��p-���Ὸ�퓆q�p��hP��{b�W�d�n��Y����Pl3IC��.�c�o��C��R]�B}�	j`�>��y����/CiV�m虪�H�X��{$�A�H�6������� �a�Oj�~���Q2���� S����CH�+��%��4����V��(�t1��itN����GW bQ�i���W;=$�v�횚�
ܫ<����+�~`��RE>k�+Y��J�ټ�'|���U���}27�m��nq$w���^1:p�n����͔����R��-����V�D�]��!X��n��%�߈^�j�/ek�z�Jq�=�wy�1i��Ѯ�M��ݞ���^�b�����o��^��G�t
���%t���&�t�BM�
��Vy%<��/�u�/�Kc����1�� y���J�P��U�St�I�k�[�iqKqq�?�p����r��)�>��)�eW=��{�u�y�%N�`��L+zESx�kzX	�J�/����t�5*!.D}�z�*Ү��� |�O�:��C����m��ՐunK�h q�g��Gd4�ZO*�tu�6��$����r�8�a��pvj��F��H�=�V�Dㄉ��4���g�Z�[NP�$0坬$�̣�H1�/��� ��	�p8�pS�7�a+��E���f6���2Ʊ��D�-~)S��jz���W/e��%<��"��(�F�u�e�CS<��"��r�J���-��ơ�V>�' �ʆ)Z�}4T���zᣇ��|��fس:��8�"F�N�	��K���@ܑ�d�RU �BVFi�Q���ҍMc�P�9="���1�ڢ_���=Y�|OB��F��%~�*qUQ`/đk�c��럞j>N�'���2�x���S��mii�9[�eGʭ��'%�l�}��G
����P[AP��W����J�SYŤ4�����O���Ϻ�w�+vv��:��g�2�B���z�̉ ��)jl�����->�ղ��zs6'�����ӯń�rBUU��H$�H��`Eu=�%�����\o��i,Z*tv�۪��"]��S-�6!��Z��w�L_��ɖ6N�Z�'�6����)sP��%�`(�ޥ��%����d~�x��WN�J[�W0���_-���/�J�o��0q���"�Ip�=���g��a��Sq�������[���]y�o�w�C�<�m�Cc�^�tI]Ck����n8]/�ahR�`;Oz]�yIdxs����LO_*,%�����q*:��� $�����Mέ��'�� d=B!���:�V9(�M������Q��Jw�%{�h�ȇd���ڹ�ޮP�"6^Gr�������L6	�^�����e���h�!G^ωE.�㢕��W"k쯿;��8�^�rS��t��ﯨ
(��="�[nm�2��	�>5BREm�}���nft>�6gD�o���Z6�m�&�D-��KԦ*�u���E�����Q.��șo�Qݻ����+s����&����ɤ"���jC�Ja����b0ӄ�Ž����9�l��+���Gw�0[%� �tlj�i(A�Y-�\""�y.�Q���H<�!�`�=�\�|H�2�Pm�ϥ�^3����p��.�G��1�$�c��ʦ�·��_)�t�`��P��-E ������t�WA#bO�9>.^]�ښ�b5A���<#�4����-���>
N��w�Q4�-`��B&~�$�)�����װ��uZ��_�Τe�0�����ğ�m�R�I���D�{h$��O�w�>�B�ȉ��zK�}R��� 9�!4Ⱥův�N�-�/M��}��o�u�ٍ�)�f��*�CҮ��.��˫�v��вJ��7��;��q�%������Aq�7Z_��I����p�
 
a@���e6��O��(s�o�P�n�ܤ�����l*5��g��j����8��<�诛�G�b��f
�ԡ�^^:�'z�׌�;pzw^��hN����6�K(1�dA�O7��x؈�NZ7�ż��B���z�S�w����N�j�H<m��∕��k~1sZ��T`N�ZoZ;�G�^]͘�i�q���E6�_���sf���l{��	R��Y�C������]�Q�N�qK5�L�|CH��T��1�W��S�氰�o�C����ۘo��~8�*Vpuqw�s�aĽ�n�T]jf�&�%�bߏf���iRϫE�k}�md@�d�1��Yd�Wr���쓆`��	۷ɕ�j� �L%���ȕ.̖�MCe�t	��y�%�5���i��i1�h�0���F��9�K9�x��2�^7��ݽ��X��;d�<,>waVfLC��>�s�;�S�2��4'섨��X	�V�o� ˊ?=�AZX_m�4[L�o�.' �o؂�:A���]=���'GGQ�x���I��6P~��_ڂ�&@� �U1h�fzΙ�S�}���t���b!� ��N/򚀿�j��%�	�I��I@wm1�>o����!>#tR+>:���4�7R����9� y/��k�HQ��6@��˳�ye�Ow,%��
4�~��%����0^_� /�Y��,�/��������T���u�v��ۼG�\���fDz��2�KY�}&����e�4+�X	S�}M\��cc���-*���Ħ��Y,+]��'O�T,�p��&�u�>"���ecZ�;��2V��F��#s	�ta_�_���q艛�<7?��WU�^Y[#D@����Ll�q�(���E�ƽB�lozDG�O�|1:�FxzL���������2F0��_K��#���$>��3k('Ҕ��U!>���41�A\�i��.������5��
���_E �y��W&)�.e��=:c��F�yJ�$��}7I48�B�H�Og���y_�(mM�6;错*SN�ͬ��0��t����'v��q3��c�
\?��}�`�e���0�1(��vT��bO��$�7�H&��F��0��Y�r�U�<�y����<e������������Y��F�w%���5 ��ם]���*��W���&3����4diu1$V�񺕳;��WV vЫ���;�.�!������9A%s�ƔB#��� �5.W����51��3��#"�y�����|����v���*_S�/Tί��\J�����spx�M�}~��v����<�'jT�*�.k�Y�p:��1�h�v��k�wy�m������X�d�u���j�.E\���x���J}�#稢>�8]5A�X$��_Θ�i���,��-�-����y4�m��� Vi��Ţ�b���4���R�������6O��bXd������A�]�I�0�-���z#4��.�tw��r��wo �J�m95���p!=�	eO�~\��R�Y;',�\iҶ踭ۗJ\�'4���Z
�îxj�Y�G����6��9�Y5�Hm|UH�l���H}#]G2sqJ�S��F���=yn�������9�aQ�3�|��Q �b���	������&���-I�c�@C�eMJ#�%��~�S��T�����c;4�cj�F7N1��3�e?�w]�Ӻ�0����