XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y9	�֎/=gC��'�����l����1���ɜN�"9�n`m���|M�x�?9�%_ȴ5��R▩W�/,�ټ~}0�W���Ue�s(�݇% ]�<�릡��g+�{J�+��<���Ͳ�����]��?|~^,c����ss�IyViG��P���4�I'�oQ�q�s�dZὰ<�Z!
h#Ǽ�E����n����Țs����ˉ3r4�W�I��X�V��Ο�JoPҾ����)��9p=�6���לޙ\I'�u�����@Vw��~�a��h��J,]�A+X`%�ޏ���)�x�]wV[AX'*)����S�C�o1Hh:	Io��5���0�&��ٍ�D!��-F��n (W�A4q���I��*AMF��G7ҝ-��N@3]�H"�?���O���0ܯ�<�E��u?�O�k���{a��n�0�Ib7^��X:�]�����ݙ��H�$0�Y�M��"�P4��j,>[��,�UK��(���%���T��U-T#V�1 ��՚�V>�^N�W�飿��O�������Ƅ�9lGV�5�(+�
��Į7��	�h�<�>ce�0��9�_$�~u-?�y�)�k���јp�:���/F��e��-~�
8�|�;E�A�����g����6����}�����_�X"P����l{#�]��)ɵ`2�<2��i}Z!��Bꕣ�V�-�|��-�t6ʫ�8],���"�.��q}\�9e�{xno�F�q��	�ww������=XlxVHYEB    1427     840?����!�i�z2"(uXr��bֈ�2�q������Z��J�N2�u�p���®����U�%l(��o��"��T��h�ʉ���iD�3P+�Q���P�7%� �_Q\�{AP҉�h�A���Q�h�Y����̈́t��VЬ���L����렪��#23G�#��6j0��'�#�beK��=խ����2�I;u���ۿB{�=�l[ԗ�E��� �+�2��퀥A.h���E]u�jH�ck+4��3��y~��������]��y�ӧ��Fq5�sN�RF� ^�������;��u����"���D���Ʉ��%��'Y4��NU�|#�[��rr+,O�%��e���KA���C_��c:S��S���]_08E gܫy�d�ܩ���8pK����Ѧ^�R���&�m՟:�#Zk"��Y[�,�����9'��ݸ0	�#��iƏ�7r�D͞@��3!��R.��I�ˮN�e����R�|.���Χe֮���v�P����y�PT��6`J�=B��S90Q,��K���7)	����U���E��~�}�z�sQA�wd}�@��L�Į�G��6_�ġ���������(P�c��ޔ.�f�cy"��Ԯ��Z���*���,g���?q芷B�MU����b�h40�݃���d%����^p긔(Sa�=����UZ�������{j�z1�`��A�J�������ҡШh�(s�~'�!��'�5�苤_�gff}�Y�h�Ӥ�w�!�����m1���}���t�z�g̞-��U�@"��#��3}�<�d��lc�>nhU]V�J�]��|Q���.�&�.���㥗uM�l��� �� Ł�cbqar<oK�Iͷ��I�.��XVD,W;�SƜ+^	��p��04ړ��'I�V�񭩓�g�x�&�<N~~)Kb}�)��,���{L��!}�#� Ԋ��
��i+����Z=#3����!V~NT���)���=,b�R�v�æi.���B��,�*�e��(ᴵ-��Am/���^�es��!�Fdz�n�w{@s)�Řϲqa(v.~��/�$=���䧈{��o9?FE��t�J�KSZmҢR.d��_Z�%6,nl�AƲ(��ˍ;���0���'��~��!H�qA�P{ �u��7hzG��)�k�����u�����3�������Ъx*�{h�!��C��4��}�8e`T���J�}��_�^Ж���L�tCQ9y�;'g��?�!:Z�y��=O��m�L��e�<z�h��Y�?���f��?r��E}j2�ukr,a�<��抿�_$�ڣ����A!�0����E�4���8G��wo�aaԾ�Ewl����V��	�K�0�av�եWf!d`��@c��F�D�^�Y�9��$���k����c�dqBȦ��2�見O�2]��yi�+��¥͸��}(�;�8��ȧ����|�Q�hυ�+��u�֓
c�񗎣�؋�Q�w�\9_�1=�"�gP"�:Ʀ>jtZ���:iK��� "�ˇ$��į�f�4������]�M!��k����IkC�cL;����ʿNO�W^c�U�x�=d�eCm=����="ax�1#���Q-
2��t��2<nY���L
/R���&��������uOS����F�rZ0��>u���5�F��Z�����Æ��s��E?�hV���/Y�,+Gom���ǚ8~<�I^*�{4+�����W�;�b��py����6�^|����!�Q
�����ӎ�vޭS����o=^�qy���ק^��U�6F2�+��:J�o<�i!xr��.B�Z�X�<�����T�>͚�߶�|�˚��wҷ�@����Yn}d��O�s���+60�����ْh'==��g�n��NƩ;8:�-�XS�Ndi �1,�k.Ə유��-��s�Lxz�Y��o���2�jsPPo�za��)>��K��G�0Y�&O�/�4˛�������f��S �Zf�<e�M=t�wP��[�
�51�7j9i�Pت�{�<a�`{�