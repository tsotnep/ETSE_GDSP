XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d�?�<0�Jr��v�[I��J�u���!2Ķ�c4@vww���Ӧ��Ku����Rm�-���%m:;��6O���"7AEY��A��o������uĽ�@��o�T8Խ*,p+��R%ʺݭ^���\x6�UŒ��]uAI��U���1���ݘQ�$�y�����f�.<:$O��0_]��RM'6��|� �j�2,�%Զ���-ɱ�I���1���/D���޻�'A7(0�@�([�d�ٙa&��.�q��ֶO%�(s�����AE�!��iD���Aa6�򫜪s����
�.�o�	ϑ�ì<�-٨,��8Y�u�	�*�)Ӄ`�w���h�X��djM���s|�����#����տ����$tJv��~�����x:E�ʸζP�]N�7���� �\#��R���=W�b݊�.?�Jh��%Q�y��ǘE�^t�wte.ʉ�[ՙ鼫4����M���4-�xf�q�I}V�x,o=x�����Wԅ�?�;'���7���!��M�������I�j?�yҙ!E25����%�.<��
$�����
��嬐�⢆��Mm�ߦc�.A����ɥ}���(֤P��|l�WTJ��]Ξ��#�/�h��
k��S)31?����LW�;
��2.DS1��&I��yL�YH`i�L�����i �����ˇ:�C�t۽+���	<!�n�l'mӎ9������x��6��7.��xcP)\�Uve��Mcվ�����Lw�3XlxVHYEB    3504     cb08��v��U3��-��OOj!O�ť6�܀����9�	7\w斤���K~79�dZT��Q�F¤p�b��>]�.>�'h�/�ڑ[���ު7�Xz���ɛ���3�U��(�ő���|D4����p���9iYf�{#�!�ʥs;����6���Fj�E/A雌؟s}LC�H�7GD��y�[rs�K?4o�0��$�I�q����ˑ��K m^C����t��@�?�1�s�s�C�B�k�D����r_zơY�x�5ڍL¦����~`灯�(����9�����q[uN��<�p.hz-4����y�U�L-u�'>��g�Ty����Qv��+���q���'k{k&7OQ���0/�\����`a�E��z;�����ᑏdY?p���旛E���*c����T�}�Q��?tuFssAAv�I����ja����?���`�Ů��s1��7~�N�^�~��%$����7!�BqDG�I�7�ےɺ�)��uB��<��pD�Ʒ��W~���ɩ�����@�z��X`.�}ɳ&�\�X$i��8���o3rv�c#�	/�a��G����P���AMQ!���?q��4}j�\�����˳DeQJ̓�.����L0q-������`���i���G�	d��ÕCR�Ӥ�w���Je� r��)�5 �3�U~'RP̪��a-:X30a�C�
�^��>�������~���.���J]�~���O�7W�r$�}�ʻ߶�Ctv�+q����W��D�?�#��!vHf>$����i��ы2%y��5�b�^S7������CE��i?C��y�1v��I�,�������0��5��$zØ��r�һ�@��;mK:�Фrb�p M<�Y���gp�����ACq�9*t�]|
�D/2���O@իK?�a�>�R��8��h��ye$��z��?����I�|�����+b��TO�3�ݠ�x�Օ�aЃ(W�����}�/|��6�w~����I#�8���e�N������S��K�%y���C��E^������s���Ր=)�O��xs���Q�Se�=����R�⛜��E;"��,Nm"�ν�`޵��âSsCoD9��T�.� �n��Z��#����6h=L�e`?��4"3�5�����I���PB%ٕ��	8�E��_H��c��]���೿uC#�u����uȤ�yX��zk�X�rK	�J����FSE5-��y����$܉C�d3��U�C$�S}8����n	�W��yYV`��׾,9��s�@߇��x��!z�WR,ϴ;�b�Is�RҺB$��u���\/A@��qH�' ���� t�9��zBy8M}sԾmؖ�nʞ�}l�����7���#��
\�+�o���$����Q��S�W�j�,��&��XǮMLNa)%��\O�0��#�۟v�R�ұ���Z��]�r�2������WQ��^��g� 
�����f_"�)�����RY��?�xG!`8kC��_�n����L2V�`8-J����!��F�YLe:^쐡�fDd�+l�T�0�S0qQb�&H\(���k%e��!.W��`!�wQ�_�/����h��61c�b�QO� t-�ҭ�wF�O��(�Ɔ�N,�<*���l�)/��q`�5�;k�P�7�7�E�����{v�[�yŹ6�i�J�i�^8���eL�%��L~X��%���b���\Q�鷀Z1��j���GZ��H�R���,�b��σn{�/;>��u|{X�;�+���e�>��b�d8�B_�'l���������J���o��	��0f��Va������?D{���a'�^��ӝ-�Zj�:� ���	LM�U���Ɠ1�(����%��W ��m�K� �7�����%4�pu���b��Rm�W�/�K��?����:�f$|�\r�^c�Gy�>���Q|g&�����H�Z�d�\v�g<�A���ƺ+-C�n!I��T�Ar{�
���p�����^���� 23a��G�e@�]C#��FO��j���*��	C��@I��j 	W�l����ֹ�]-��t}�s�%}�s)Yd�qn�-{$5��b�'���l'�;�5�����2X.�)�7|r�3��r���P�?H�mAk�F�(���^�&V+��E�fb���̒[�8'��Z��/\�y�ϟe%�����x����
V�zx�����8g�����M�l˙P\�Ki�
?�)�0��$�]E���~L�b�;�{!>�������;X�	�Lt�7yU���h`4V�s�o�o��;�3�b��mi����I��;2g����9:J��3�αu ���	���:��/v�T�ã������{�Ʉ�<P�-��TŇ��098�Kd�(v�g�C����X��+�"�#�E����u�e�73c��cu^����4_p�D���>��!�-�I���V8�6 b�'�K(��/�C%��â�D�9zL;Z�/z��ق{�Ja}כ�C7Ԧ��)N����1�WP�V5&Z��5�/ϡ�D�r/)��} p�`��M�Ę)��.��!�	��판t:�U�QIN�ۇ�+���r;G�u��L*��e�?��r�nbt�ϣ1ohB���KYrĤ�T*�ujH�t�W��� �{�(�M�Z�&
����FBG}C
?�s�^lCy�.��m���{l�T�1��d($i����8�������kR�u�����lH[��D(��MBN��rU���,��N������������I^�Q��iM�0F�T$/KK���G ��ƸPvOc�-;��8�GQ�a� �Ё/0��/gw�c�z��[[T]'���b6oO׃��%�YW�B��0���H:T"Ȓ$k썄{�M�v�yp��������un֔N�=�{u���0)h#:�&����PW��"@lЪRA./����(V��%����K{5���\-i|B<�(��hG0��2�*ulg,��$I�aP���t�=�J�Wu�$�ԁ4Cc Db9��~l{[����m(4���a��s��
2���c~��]�PZ�����K�WK�w�K2����t�?Q�*��t)d��G�z�R`��p��NO���r�p�R
��>q���!Yc����\�ￇU�#���d����{8�6Ù!�˒���������R�G��