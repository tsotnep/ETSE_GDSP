XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�Dڌg	y�+�0�"};%�Lz/q��v�;�l&�_唻��	yE>
*�YгA,=�f[����H����@�L�x΃~��\� 
2�M��_Y��#��>3�S���xW|M����� ?Ѣ32���
6���uu�k���*Ozl�ǯ0\�-�\K���7�9����=�'�a_5���}!��5W	�`�]��;�.Yq󄲩��m���J5|�[e�`�3��E���7�_�n�5�t	�����o6�W�i� c�C��g�HFĞ�1a��f�]_P��p�#���@eU����b�J�I�Z�_U��SB'F���Ŵ!�ڶW�|	����k!��Q����Ũ��k5 bj
ݑ�=��X�����3����L��'����.��_�?u����"���V���Ӡ
&�6ST�=懢R�"������Y�l�1답�fz��Nc~��7��z�d�(���Q����*��{�ǏFӦ�E�>� m2�[�L!��cH�J�?���
`�\��Lɱ�r���v�^l��%`V4�	�+���G�JP�)������ʸ8�GK�۱�!�v�
s#�7�*ͣ�k�)!���6M�m�E3��a�݀��xE�i�'�F4@87�r����&�ܪ֎�D�%#���ԛ�~ָ0x߽���,�Zہ�ږL��c#BYG�D[nC��5Z�Ə�H��8{D��{���(* G��z�Kܫ<A_�o䓀Z�-�!��z�C-y����y���˕�����+O8l�88:XlxVHYEB    fa00    2560j�Ǿ9�DEd����'o����In�hB�tdm�,��81����n9��"��)53H#�ad_�h�݇`_���D&�巐A�c�����eVwv)�ϙ �K��B6��twY4�{��!/�o$^g�E<���]�"����wO�|�@t� бq����� q!eT�Tiic%�]J[�������R��-�Ɵ���hTd�(s�f\����!��[uYg�_P����c�7'3eM�[aU']�f���q!��'�@��c�ؚ��s"�?�l3�ҜbkjD����tx��A��fD�9^���Q���S�8UB�'��E|�b��p�ܭ��t�ŝF�#���N9���6X�
s��*�&�e�i��ڭt ���jI�+HY�����뾈9�G�u�	.�=�t�$>�(w��$0��BϖhCmN�'�0���3�l�H}H�xHk�j;���շ���Zu(I�0��Wv�>�v���%��"$_�x�xNƌK��g&����E�FoZ�4��g�C}[ޫ��SiG��kf
W� ���E�&���|)���g����d����Ρ5��t����r���y���NܽY/Zi!��mÏʁp��m+ng�XvUԂ�!~�^NG^��4oUq���G���]�y%���Կ-Q۴l��N��;qU%������5F1š[�Ggu/����I3������=��:��D���&��O�}U�*�=�Q�ݮsȷC�0�݁4a�J[�-�H������?��BfM�;Ej�Ղ��c�|֘4|��~ԛ�uc�.�0���ǃ�6Y�9��D*�a9v�dl���e-ZM��|N�������t Fc����%�(�p7�ܺԙ�_]~�;L.O4�b�.���0_ǉ�1�]�ZS�`�i�H3}�tې�b8*"q$P����I�⛌O�5 �0������%�3��JƮP�!���� 㔝�����X�Xe�8��Y`d:>λ���Xg���¢�(�,ɟ�\��v��0B �K���;��7��ߟ��7����PS_l���J���H�����؇r���z��i{l����inʏ�^zյ�2M6���g�;KV���Jz5�[�S�"����6���D�U0Xx�A�k!��i��:�V�	�K�] ����D�
�:�^��u�酱}I���3��L���<�L��Q
��������;v�W�-N�m%���vA��c�m� �.�tF�FXBY�kZ��<��&�����Mm�tc"@s�@ʼ���X6�U !؆d�!���^*Q���*o�j+c��������,4{�BX�kc�<��{p�h�g��U����ᢝj�ϘB"�D]���k�&"��-謇U��|�d\ܠ�gULg^��E�C
+�g��Rs�KiE���BJ���a}��?��9�Z��G�)ZT����z��/�X.�٪�5�5ش$e�͋�n�)��q�t�sg9�$�Ii�E��`���>3�}C°�v?Kܞ
�3Σy�����%��[�'�+��!����`M�������T�Gf�RM��Z�usO0�jc��>h�C)`�</K5����9VLm��Jr��sr3<���#��"\N��@�N*I~(�ؓ���&s����cVзG69��B�
��B�P{N����vϟ�*�f��
�-T�{3
���8�ڃ��FX�ކ(Y{-�@��{��h?"��;G(��
��1$.�k%��h'�G�rbrԬ�%s4��F�V�� �LN�HF�e�1�E�����x�$����E=��SG�3�C�2j����+~����9��8��Ci�b[c-c����EC����-s7y����z�@�D~/��T���)�a��W͎�d�=piS�}�i�ۍ\m�9����|dv������9G�Qܟ���|�������%w;#����E掞�m�&��!��	�9�LVy��������ӛ�����7%�TG��&T�Y;z]'��"h$�{^�>����B��i7/S�@^�,��I�&��.�%�ix��0���Ea��Q���@뺲��W�����M'o�~|KU���2��:�0���z�P�v���>�$�G��R�,̰�wd�ZcG{�Mʃ]��vyJE��3,��R��I/}���� Cӳ��k��I߽5��(@�r����g�̝�<7����>�95w�ת5A"��1h
���J��^�'���7q6(d�R��=)+����/q�q�A��Z+M��ǻT��k>��D��g�,�����ڂZ̓5��J��P�q���+N&��&Je+%~s�$=s�zVo����k<��V������[Ч$Pe5�5�߰+���1颸c3,�x��mKHJ7����0� �-��P�~iQij�r�`Z�UV�Há���}�,vS�������{���`�xQ�j�X$�G	����j�;��H�DU��xW�^U�K���#������72�� ���U���Kѵ(O`�V��2��a�M�N^��{�H�#��i�ro�0��77TĄ�V��.W�ې��*--�K�sa��R�����-Đ�V�i�WjcO);��Iz�F_�L�q�mֺ�FF�e]�����[s0���2Y~v�흊#?��Ĩ�MҲ�l[e]^��~��{2���M�-_��Z��,�Ak4�m���/�ǂx~v@�ڔ6��j�cpIt䒠/��� �J��q�D����`�C��>�XëNWHKΞ�
�����c'��E.��� -j�^tfM���%��lj
]�����ۆ9��~�K�<#h��RH^K���Sq� K�<�$Ҟ�wE��50.�-&�+�����C�a�v$����8�đ��h�BZ̗��lN��_���#�������b�'e�0R���Mv��x����P���[X�
S*���ʾ��( ��{�>����d��O��w�Cx!����
k�#�Z���@O��?�/W�1$�9:��m��WcQ�i2*����M����-�f�#���%�R�ݤ:0��l~EN�=�J�VȨ�Ϟ��<=[���_Չ�=o/Dډ���`��
�f�{�u����uQ��2'mp&� %��ॽݭ4��^�%��� ���׬��yէ�^��91� �.k[f×�d�s�"�	�`�Q_��Ȟl;'4w�9�:Z�_4���@�j~�?�(~9c
a�i���D��3�s�!�,똉�x�/��O�(ZL�vW�'��9D衡����;����ո��B��ڨf��O��YucΝ~XY�#&b��c�$�k�2�2E 	�|�LX�܃ߞd�!&�\P[����N�ϓ��l:�:��к u!2oi|�bC�N
��` �	�>`I1T�f��j�y�͝�V�����Oܒl��A!n�|�2�	���//����ǌ�A�v�naxƦ]����Mо�_��J���1�����D�S,�-�zb��%��u���,E�l�ޟ�6'��S:���k5�����Ě����]�8�BS�ܝu�e��8���H����S���	j�W�=��"���t�S�@7��+\t WS֫�S�7%����q��߾]U����W9�1�g��s쿤�m}��~��Eo�6tn$���m>�#L��|�֔"�7&����	�5&�x��WZ�_t�j����������=OF�a�ۡg����|9��6Lk��F}`�9:�C��=y�%���U��%=�ק�\&,1�z�hU����~dr�L*Ʀ�ε�{̢6��V*����
�Ǟ���!%A������͠,9��`N޼�W�4�k'#R�Ec-�c�[Y�ct1r��Ғ�a�]�����=7��¥_p��[[�Pi��HCSQ�������t�.�z�Nj���>�F���2�딎)5�����}��1�W��-H<��c�2!�5P$	Xs�8�aR�~��`��3�9��{3fn����h��kn�rm'-��7:(�ؔrF��;9�ݲ<=!پ0^��l}��LE��ց����W�^�S$��L�}|h�|sO�g�$��ޜ/�$
;`�&�l�������pݳk�/h�\��f65��!��ND�}}aŔ�'��N�<��_���SB3�Jµ���XR:3ٜ�����'z��M��s�'�������Ƌ��_=��w������?%bv<۱w&�r�C�.0�Y�Pk� Q��Aơ�j����F�6o��8���qbk��=;y9��Qj�8��'A*0����sI.�b���r��R@�w�)ˉ��n�#mż��◕�{d#�t2;�H�7�CK���*������ �0s@��W��$�~5���z	"H�1��F3�X�]TH���6��^lx4�r��؆��z��/�Z�?X�S�A#�_�0�0�7l2��i}PJ�p�.���J��e��V�3,��V��|���-���E��?��>�M/2;�|n�qзՈ����זJD�-�+�J�j�]��M!MX���&�(BI����V?�_�.]����^y�7�RAMj� �[�������Y� 	���;<�����6$�[)XKJr>�[�4�O�EU��x�����-����t�����ŇG�����m��)�꼷\��do�����wɺ}�V�;�)��F��'#ge�-x8>�.� 	L�h��H�b��U������c�r�v�o3�`r�����9�ɑf���;����)�=|�������V b��|Xp��:,y�u�o��]Y{����AS��-��$#�/��CCf��k�YlJ%
82��H�[Ї�0�HŹ'4e���6�+�9�7>��b��$���������[����$���>쒐�c�9�"Q�g	���t��ndZ̖2� ^���>�Hh�;��̪�/��nY��#>�KF)�סCw�nQ�%���Z�#�N��_a Pp_�6�*F�Iiٜ�<
��6�΃�/�,y�ym�zroͭ�[=
�x@�R��췯��)����+�	�j����X�	���2Q�
�ҷ�ç��t����G�L{�z�J�2S�X#ķyإ%�}� �L���H�x���"z��edj�.���$L⦖����v����5*�9��B�,��e��BmB��_��)���"�4d�}v�i�B�+��ӻ�v?O_��ɹ�+��饼I���?�,�Xk����w�O�������K��s��ѩ�iK5 �s.0���u_A�|���ݴ�^���sW� Q�f^m`�֏w��j��=H6-���'��5�cg������������������ȱc�0��ű��^�9�'\���ı����>\�ê�~a>�$6�!$C�N�&ө�����e*�x��T��5Ƅ8�e��Kl��f�K��߈@�,L;o_	��&�b��CW���;4��s��=��<"���Qn��㥯�>�ͥ����9��E��kJ�c���%��	�;��Wڌ��T{�r���.7��.$�̓Cp����/ q�TKS�Vy�����D;��=�jOl���_$�:��VD���R�.g>��L�	bK�o~r�J?�2%G���O�Ӳ���� /W�f��咝�	�>�jַ٢~��-z\%o+�����M��_��Ъw�.W��=�{2!��(���}�"���(���
�ϱ��s* 6˩2_�ږ�7�H�i���[�*N���~���|�奛iV�6%<����:¶(�ס}��.t��4�eR�p����Ӓ����^f�9��~����tR-�,ȴ/c1�=u���-��u��XB,�+��u�:D<��5��<�"8g"05f����j=l����n
���&��W!��k�"o%�o�R��V7,<O�zt�l\�)9��~��ku0�hhR�xĨ觺�ZW�S|Y�i��,�=9�x�*������eB�\��$�Ic�ط,�N��i	W�����^��l�5�ƚRc57��&'�2"�y�*����e�K��4���X�a����G  ��Ӳ�VP�L��d��3�L��RT�-ͬ|�����$!{
�͜sl��7H���c�[ �8�z�p����vT(��O�s��r��6}���4��е)7�DY���e�f�]�Q�̸�*���BiՐ(��.��$��sj�� %�!!g�8 ��j(��:d����:��J��@"�F'5�ƣ�LȮ�{�Q��ֿ�5�	SMdF �DFӰ��J���c�\j>�aA��fI;ev��y? �=�OwWMǒ-[��}��K\^�����NA8��߀סYہᩫ�p��鱘�����)U��<G\�UQU�#�eY��r�4���h6v�u~�����O�7�7�%�┛��J�K�b��A�PϾ���\!�zd$��`20Ee޷��P����Ɗ˝�D"��l�Lv����x�3���\W-?ڔ�O�c�{��������Y{$�z���󬇼�Ù�%}��C��9>ϵsX��U:V�|ɶ7��Y����Wr}Zg�|e�tLg��J�蓑��l�#�o�ZosN �܏��|��w�_
֌+<Fm������W`9�1 㞣���1Ңp~�#lɊ~�]8E
�21��6�Ǘ�}U�ҽU���y�k�-���f?�h5kJKߓ�/����u�W�w{�Y���1�g��p���=i���^�&s��Ӈ;85-��I���SC����Bh�b�V���ZL�*��XIq�5����*�"ޢ�'w��F{���E�H����2W�f'B,�X��WUq�S�v�Fʝ4kp�P�͆�W��K����!u��߈el����C���n,U��D)�����[^�H�N�C��.\7V��_H���N�"�� Z]�҉��Յ�6�i(M#P�$�&>*N@b��ڥ�n����T�e��<�z2�n5��@T� ��D&�g*H�VZ���Fg�U����:��vn�ɡ2k�&m�J(ĵ��D�@��$�,f���r�3䁖�{��<�yS)I���BTM���5q���/��"�#�̠�k�)�O�ɕ$Qh3f!C_XLi�˥e|Ny��@�aI���M��8���l~/�s�&�{~�[���`� � (�4(l������R����UWj��;���H�sL�#s̜���ߑ ���>g7^���h���N5B��I�HG�ejg�h��e+}�f����1ҪY3ӄ=q�>�]�TZ>�9b�a6(�sLᲖ�a^�1\��H���88]�6�//?V�����W�Q��dp2�H�����U����	�v��U��@L�<\p��A@ko��G�H��4GQ�ؕ8�Ek��^C�'j�D=j��<�>Nq�x�<��l-�2�w������wp;�5�O9��7������F���ɔ)Z�E�a�Cz]ߡ`q|�H`�7Aa���~�Z���=�.��q����#iL�}y�?�?3�`�;8���E��^>��g�<B?��^���]�Ҷ;&i^;K�V/�4\�?=9��/���0A��[tu�|e&�S�x���=t��{�F_�" 'vF������-L�Z'�Иy��aS�1;Nuo�F�՟b����H5;2'1cL�Y�g�
�R_�7�򆐺�D�rק�}���h&_�d�
�eCr)�?-������-�"%�2�rO�h&"�+�ɫ:��j{9l�+c������4�W�D����(Л@�V����o$&@�Ji)D_�f�zLgX-�ߛ�B&#$�2��lP����{�y�
^�<���b�-���d�������8ĩ9t��&�`�FG��x�ػB 8��1 �m��B@̃Nٸ��p�4�pJf��%��H�I���B���k�fJ�p������Ti�
3���q.cg��C��
6s�Ő3��	ؿ�]6��ѿ�%� ��p(jv���Eޫ���k+���Rd>qL����eKf���b�hF��ǰ�`ѱ;.�!�i�g�u�A�16'�ه80�T�p8�\x�>�˫}��4����������o�|{ԉ���<���8A��1w���s�==����3�)AX��j������H�k�%����0*���3���{���t��<���l���ꞟn?"aa,kyyg"1Le�>25&�ا�j�%2���O	�݀��$-͔��]�������X:���A�.p�����9 �G�H��,�r��9_��G��L�޺�:�L��f�.��h5���ä�1�z鳩�<Y7���l��j7��(C]l9F�l�֓�_Bz'Z�{�'5դ�<���mkzVF��g�N�1qL��6���+mS�P�Z8�ɞ��#�S3�J�M�Q,� )B�9�U
�͞��[�ӟʴ��o��őHO���P"����*�,��5��\~Ć�I�r0���D�B�{k�ՒZ&W`�|�������$A�#^c;S��{QL�2���+_p'!��|�%i⁃�TG�=��"S���0���w��APp�J��\������D���ˣ�?�=��.��"��"GúL'̱�Re"�`O�n��i���(	R#�wp]s����;Fx6�b�x�m�EK���$�Cw�g�����uΝ 
�	�B�oF���lj4X<�����(j���e<̪��tBƨ7to��^��㧃L�/
���R���#~��f�z"�)�Rn�`Ș��و<ny)o�Cr�l!Q�����'M�-�~	"!�7
�P�~wk>�� �4�ٓ_�4�t��,��ᖗ�cj��u�����af�8�bL+����ц�a�c]fv1�^�w pRc5�#�%f����qr|R�d�v�j�����^����S��zĚg�>�	��~��%�o�1JiR�x��/y�z�Ye�����DG�,��mn�O�i����U�����!��?�o��۽r Wŏ�{&��ay�Q�.�bt�S�-��0"�$!0R�^1k~	���+��;��������0E�C����c���)�ݐ)��'����֦mf��]���mRm�I-�zV�Tlxv%.��a7�?:(LT	�
�zg)Z�&w�s�Imc ԕ��e��8� �-��ED����IURJhxЦӪ`�:xN)���w%vlDS��W;�~�hm�
��/���&Z�=��Y��-�ޮ/j�<qb�ZvV<�f���aW}W���lp>��d���Hpc��l6?A^���B�j���/�K$ŁP;�Cs.,�� t��"���A���#����Ա�����
��-�(���&��l��䊵�$G��S��Y��A%�X���1W�������&�t��@2.)^�{�Q��'��J��j%rG�x��V^{�+	����("�ڬ��)�ӽ�ۊ��z�X�<T�XlxVHYEB    fa00    14b0�t��`@[ևa�<�9�]r��P䠙瘢��2�U;3_0t���>y��T�8	6T��u��FS��֤�( L������i�S�g<z9\[&���(�
����Ē<��}Z0x�蜉�$��E���zf�E��` X͒w��Bx����mp����V�is0 �ĺ&���:�������*��s3��v?�>7�=ϕ�-"y����wܔy�D�
��{��:�VT����p�q�[��tzO�W�XB;�.�/|�N�}s��Q�t3i��=���į)/�f4��T1<	l�$⪗I���;�%^�H�����bVIÌ}Ʒ�/��<�p���{��P˅N�}F��v����Ed���.��bd�]\�g[z[����h�!aT7 4�'�RМ@�.��M����+���6C/xx��1�PU/�a���f��<2�7�R��*m��wM	
B���b�C�p��J1�c�^����gy'��̈I�����1Z��� <�s骤�'\�-�&�V�V:�W4���UD�D4R7Ot'�n������&%u;x˙v��6笧�]^MB�6D�[|���Ċ1��vi'V-a@��'v��B ��K�)��\�z��T,X�X�z�+y,oL�6A��-"��`b��\�5��V�O����	6��%A�����p�^�f%����)W�Y/�_A�
����OZ�߆�<(��o�,5b��@���H�n�xy�5%��)�p��Q��|U�U+��N��B,V�[0�`�?���jj7�h\��y�kzN?fqe�ٍN�đ�HxB�u�\�W�"�ϧu��ȗ��Q1���6����t�� O�"�Zb��.��P�����Iәm�v��\��>o6ʲ�B���Y��}r�%u�;�[7�:(�t��3yÂ^N��\cm
��؏;�*���]�Z0���"��<��_���bsޅ@��de�d�:vdaQ�
1�r����q3Rn�n˞���f�����NE=�n�V���4���V����u���>Wc3�o�oգaA�]6(6_JM�۩���� �5
1�٠0�#�s���"�	A<��m���7��6J�t�H��5�?R���CDx��{]���u�7&cP�o��i�a�hj��/i>8���>bt���9 I
��d�&�P���xMm���l�Ly���&�M�b�HK�TEgW��[A����`�H�汿ۙ*�G. 
��$ڹ'}��
��jD@!�B�`��-Q�7���4���
�6M~����K��r'�O�"u)�K�\%�� ^zD��>���"1Z�z��I�AN���?s�	��"!5w���}�}��(h.#em�g{���F�W�F����z��o�w����R@����J�X[}���N��d�㡿�$Kn@#C�}{�HC�͆E4F����G'�k�%]T�iE뼕g!�6[Ɓ�B�-H��%�Vj�b~�7�BT�G��ZE6��W���f�]}O�Q�/�̰
��ɶM�B���c~mZ��<�xwfM"�0�[��� �JF���j�@��o1Y�Rx��Ju�A�25W����T�,�Y��Fx���I�����ŵ-SHiY��-SZ��j�L���'Ś`;Ufr8�W����7{��AN�JĳF�;���X
_o(R��-�2��~ �HKN�nM�SF@�?��T+v5�g�rϒ�מ��{��}t��`x�d}�ԱoX0`�2c����.�Yk>�N���:����9!�p�1 �IYe]�3��M:�Dn/��u�Ӷ7|�^��ւ�U�iS��.��M7�PV�⠱�'�-8�OGV~x��2̇�on��
�e�.�=�QX^=o��u�7a.�i��`�ύL���f�	jr1e�����;&Hb����(��ub��)U�LN�F,y��I�����]X�7��sg<4�R��h*\_��6���,x:
LbX�Դ�B�'�E�M4A=�q���������hׁ��o1z�?2~�*R���-m 0\2s�)�Q�ឺ�呠�kGv4R��G�4�����<��������#v�`�����Z��Q�˄tmZf[���(oJ��/YA�U�l��`8�(b�+�I�\o�D?�T���L�?K�������{���G|�ݒ�#(�]�iU]�g�?��NLU�950{P�%b���lD��6EV�jWփ��xퟩ�H��'/A�3$��+,T��ӓX���Ő9M��YKy������h#�S:4��@���$������I�.u�㎚��:���Ś}���wI0EN<�z#��o�9��998[���*�r]�G>_Ć$۸�+[�0u��^.��[[�"˃=�=�W����p9�9jmOC}��j"Qy��O���}Q(���ЮBcW�R�&(iZȈN���\�rR�6X�Q;R��Z�FEq͌�k}��ou+j�N�(�iIƖ2ҎR#uȸ_z��g[ҵ|��/�����@&Ш����%?&y��.�z���Q�t�,(�D�|��	e���i����8���q%���}���Yo
�|�7�����6#�lD��uXlY�F�pXo�֨|�s������٭#403ט_ӈ�����aS���H��(�z/��ֆ�R�~���Z��Ys�ԊjB��.��I@u��4�⒗v\̦e�Z�'�5���!#Z��WD�4�u��-d��m��:Z����P�4����*�>�����5f�~; �{-���g�f�i�8ҠH$�Vp}en8,ㄣʱ6�vx�� 6$TcN�/f:���a_w�S]�ޏ�F��K�a`���F��}�y/��S�w	R$�n���^���LsO1�B�7�~�<7��}�����,N�q�3Д����~�T�P�b���x�0M��ځ�0�(��I�����Z�֡��Kݤk�_2���!�;y��82��� �RS!�- ��b��꒸�x�n��%Y������>c,�R��s��Y~����}�S�߆I��Z��v�^�����da
�ʼQ�|n�Ƶ
(��;`{�mW/t��;
U�a��o]%@�2j# ؆qD��pĸ��1R�w>ȹ�����u3����l=i"Z��j/a>�Kﭐ֜���Ôb��6J����m�#�3>��$򫝨_j��C�Nh@g�ڥ�n�~����ε�Fu��w�L=q������d5�±����m�}[�g�E��}�!�fb�P�
ѓRW������)Ć�N�xLȥ4����������C)���N|�@W��ܖ7+�|j8Y��i���OP�̚I�<F�|Ko?����������0��=�j�G(RV�5l���{����$��r�t >]�cPE�9]x�^0GdTx�ǔ+`��7�eM_J����$�w(�sm?�����WG��!�w�g_r�4Y��w�r�>���s��|:���O�u�����{���S��p��$�y�>6rok40���@�u��ӳ˾[���f�3{����T�j��ђj��%�Q�e�1���u�g�R�O!Uܸ�H?dQo���ť^��)C�F�x�£d}�ú�jj�gI����2X�C�i��*WGa9#
�7���}k��}�CF,����,9nÊ,v��2گy�����a�YF������>![�EO�C}�o�J_v��p�����Ɔ�(��c��y�c��ɿ3�V�0SЪk��[�����UG���ޓ�*N8.<�;	f�9a��~����\�g��%mOk�����5ظ����4$q�FK�Tm���%7�ix���=N�6�	wh� ��s����
^^u5WP��A{hZ.��B��	e�6}�]Q緝^YXL�j�ty�q�3�Į��KY"S�Jg�1�.��14*��`š %ޤ?ͤa�l�J���\��g��uϴ��O���/i��_��!���N����g�{e����)z�̅}ʆ�l"=����9�#A�~�@��w��R����{�|W:Q!&I�G�ki��i���v�и��e""��l�X*AVߡ"�ظ��A�,[v��-u�H�H�Wם�j�y�y˘�>Aԝ�]������o�O�k*�#^HU�>�M�=��3���k�،�_����b�o=����x�G������>b7�D��Z��'��44�m�n�oc㚦��EC�̗a�ƎzLa%�ctF�� ����C��0A	ή^8����Xcp%;�K��ڿ�y���d�_'S��O΂Q�Kډ�
�kQ�J)Le:��fRn7�K_A)�����	�U��FT���� ��c6"p��`� }_)�C�ߐ�B-�l� ��ZiJ�eĞ��:E.Ƕ��t\���Kk��&�a�镧DQk����@5V+k�ژ$a,�̈́L����v���ѥ:�mȾ��_v�}QZf$�ѬĽuP^^;��rp����E0D܁(�y�h�rR	�X
���/XMg�4fh��5���	�F�3K"��Kxץ�!���q���\ly��ػ��#�.A9B�_�ɟ�ďP��?Nԝ��_��&�.i����;��!��4��5x��t%�pJ���
e��.P�Q����B�B9S%k.g��e#I�re�x��M�5�O;��r�9���> 1J�s��C�F�X�rUP�����~"����84��`v�ޚ��S��+lű{H�S�4���X�����[�1�1��-jg;�"!�7J�6��Kߟ�	�
�~ �D���p�i����ׯ����8
��X|��4mh��xT��N��3A=s�b�߂��'�v�I'��(ZB��+�)��LX�d��0�� ˘D��0�YxU��Fʺ�N����Vv��i'1�EľNq'����eC/���Ů6�EaX�.K������J��y��d�IV�c�@2�I�!�����=�1�A����s�X��T3�pYj����!`edr)����Nʊ�kM��_Wϑ{�\Zz]]ok�&{\m�xC�������HIi.� �>b���SM����L�-Z�3����F��i��fYV��[SJ�����Z�{e��G���*0�`��I�d��z�TA$�ެ]3a�arx�v�*ޒ��T������P��,Y�+}�&T�HC�ZH��k��f���έ�b|�-��49��o�����-��LN�
٤2��Yr$��i2�5��%���n��V]�r���4�uW���@xQhM���x��O�
��l�^T��9�'W� �����\o���XlxVHYEB    fa00    18806�wH����#*��v�k�*�O)���@"��wl
���6���a+eOwB�i�QM�S�Ƒؼ�4נ�p'�8�h��(�];z^G1���w$��
Oϣb� �5�Z��{(O��q��_m� ��h:l%k:Т�n?,��°j�Â��s$4�")���s�����Ev��<���Y��z������:	�J�	:S���;x<v-�k"��kE�p�I���N����*:�b�i[L�z�1/�n�5�P�v�N�U,T��
Y�9�z�M��ew��g��"�!�&F�k���&%�L?�BN(��p&.����@�s>a�Ϣ�K��R���ث$`���b����eֻ�p�z��F&���ߟ��L+'��������f�.���:��Rw�B�s�.h ���[�� tsø�H��ܹ�D�~c08Φ�&H�۪[��M�*au#��}q���|�������T����m!�zۋ><��6	=��E�e�5/��:`�%'��(8��V�v�K�յ��H6n ���w-��t�pCyM,�۶���M�ؙ��[0G��3���2��l���m��I���"�>������Y���a�4�㴬��/��j�tq�FR��]��Ã+��\;��8TZ�[�7�
�(��3�[k��"��j�5�a�&7�;o�tAV�*�&����`�Dy$Tk#5ZN ���8�)!����=���9��������	;�߇��č�!��,ԁ��,�}2�D)��Cr3��?$m )f�Y���{^���9�n�\"c�>(R�vꅪ՟S�X	�HC�@�x� i��'UG��Ĵ�x��3���S(d������3�fp˙�4�a�qwL� �Ń�,��IK1�!޻��t^cI�m���׸M�e����v���&ܠS�Գ��� gS!זa�]a�*�q�k�`�����w�O54_�7�t��v��R�@nQ�g/ȧ�kx3;'/��|,����=�K�B�l��NW*UR�/Jߪ�l����"g¢3ru:J��]"'��g��n-5�9���a�:�ޝ*O���T{�����-34�ѻ�O���`��x�rg)�S	/HU�{�Ӆ�q������>'�N��]��uU/��_����D���0_��Y��X�Y�i�5y���n�M�8`dɵ�vk�CO�|)���U�������_e,T�`H��6%`H-)����R�f���}l�����V�ډ�F��V9 ����%���~)�AWP �tF`@?ҟ��A�F��p�W��Jf�-���M���S*�X�&S�l{l�G۠k�/�P�`�v2l1���m(Ci�Uv����O�HΠT(�uö�x��u�*���\� ���w���jFL��ޟ���s�(	��31�1C�I�L�ڎ)v�tB�tZ����	֛�8n�[�X�����6�eE�kJ+���RF��Fb딊ku0�h�ޗ�Y�
���$$)�8��I�qޭ�W�a�ѧ-�r2�ř���Ù6Sz��OF��Z��Έ"���-�{�\&���Ġ7��º���m��Z%�F��WE%�:?��q黿2j��d
U���T.`��l߰��J�����4�R\��=E π1Z�:�9�g��/���7�⧽&��ߡR�J����h���8��o��s��EX?�U�!�;���N�C#59��K�ч-|�S>��L�f�ņ���3������[�6�SP�?0�c7%=Aj�ttU��eA���_�)Y�͵x��Ժ:�;#l�d) ȹ�XU��w�Ilp,W��`��g������#m�?��_�`t�I�c����z��Y}k}�.?�]}��� \2$g&[��Q�[�Jqf�w��{�#n�����e�k�l~U�� V�\A747�u��K�ܺ�EK���Jϸ-��{VO���j%�adj�dR�o�9��g��=�^ia���o&��>�3G��l�����4)NI����XF��=x�կ�4fd[�ƕ��{�|�@/��MWn�b����N����( �TAV8/�̈́A%<���K���5�zİS�5b;��y��G�'ک$�#tⴧ�z/{p��e����Mb,:��.���z��E`�o��gѐ3���"YL4��S:l_\��R��QU���fg)K܉���ԛ�j8�q�i$�*�_��O`��1Q�)��N���aK�V��Q��:�LRE$�j�8u���A��F���cR?z�9	�}�{���,��غo
��Y{#$c�������o�������н�-z���
����L��G�)�D*�����(&��f��W�صNQ��jIX+����4�ᷦ^&�&��j8���?���� | �H���[̣���k9�g�#�Y�l�R�3�U҆=������Ӑ���}��f�=#��h��ǐ�<��an��ƀ���u��ѓ7Ksy���ud�|ڼ��A��T`�"�c��}Q����熇�����k_e��R��D#a����o��o�5!%Ye\�ա�$O�;Y� �%�0�V`UfH�|~vfo�"1鴘�i�0VIۺ:SZQ�ވ.Bm��r@=&��O~=�ǘ� 9Z�cn�ET}�_H���T�BW�N�����kI�H�M�&���wC|Ҽ��-ٱϷ����c���JћoH������Dēa�	�ɻ1������>o�����A|Pg蒾���;pC͕�UL��i������,XՋ��Np��5��,�J����p�e�Ea���ޗPʴ����/��Y��j�b��x`2�[��+N�����0@R	 ��>%g.����W�A�Q�{�@P����G�"E6?kT�Uu�ߕ���=�������������Q�a_��7|Cklm7k�E�ō��jƒ�@�v � b��2֙�k����L,�����n��L&���U�"zy3
�K��Q��ⶄch�͚�2�X��3�������4oؐ�0  ۓ�2��&_�B��+<����A�� �
����oy�)0�����n`�8�aOL5;�iQ�В��H� �]�	u��+�s��s�6*M�)6�|'璕p��f��Q�.���E
�/���K=�&R�����8���oD�F�)��16�S�/+3�Pq�D8�X������Â��˅�Ft�O��y�6̋��`�B���ϣ2������K*�|mlԆ�4��H��(7S�q ��k��A�q;�u>�%�h�?ud����Z��\�Ԝy�d�;��n��S��z!Vk��n 'G��m�k���seø�?�p�T�ݧ�4o-Y�t�83wCa��Cq{/WW}K�&g ��9�i�1|\7կ6	���[���8Bq��q�� �9��>�bg��務�`]��vųФ�8JI툌~��g�LU��7L���3��g�"��q�H�-��$NH�E��
נ�	� �X�:�6P���L�-�%u�ΈUl����b3�.�a�佝�|��%NfP�#�����ҡf\�^س�uw�T������PP��Y��~	�wUi\����P�Prx��_?q3��']�����7FFH�h���Yh#�ǒj\9o%Y1>�z;��z���
�����l�y!H���N���u��zԵ��BH��1��?
���q���#��T��3��9GAy��".�n�����ɕ� gi%�K�	�h�m��W�Ǖ� �xq��R� W2d��"A	�t��}���{T������1S�ʤc`@�P���g�������D�M'�1��@� }�;�n�\M̧FS�L���;@�b�odø �F��,�2��b|/.i��A����`\�_s[�=�Z�G�E��gQ��;`��sGRa[��<f#a��o�`�zfbt�r�9���Nr�!P^�ph��M��~�Q^^9U1����$3SU�O,r�p��usT���m�%������00�D�N�E)^-�>�(�����c���Wa��UNqcV�3�b�0���a��J�wM�S�:��7�1rkV��i<�f@`����ߢ���y��t�/?���C,�:z��XSRl���fRma�E<�;�>��%܊pgYO�[�\��lD�ɶM{�W���\����7�	�����_ҟ�-`��$�����4%�0��l@����V�P�X6��a��1f
kY�b��9��B���`>խ�~UJdqW��~���b����d.���$z��X�=v%}�d����5fY�y]��5�����6�-�;�;�C����,c"���p7=�_�|�2�fSoN`�����v���Yf��u!e�൙�I�3��<S��]d
L��V��z�DG��
��BP�}��&�W�n��OR��)Y8�ߙ�i�.~�#&���[��*$��� ����W{����Z�����콇��X-��}���&���ii遬�8L��'fOwFeNC gO�`�'����n"��s��0\Y�a��izB&O�������ذ�A���h�9��/���l>R�l{c��QpcA�I��k�]�ey�ӿ���8�k�h�Ҧ��_.�`��q�'�`���uʹ����C����s;U����߸��E~U���d�� ��Գ��@�.��M7x�Щ��%�����S�fIa�Y��l���(_���j"d|�;LM �C��n҂3�~����0��1�l�VeZ��A�I_��h��ɫ��>e���Ɲ��rT�ٿ�o�������D.3�I��NdE�m��2�ۈ�W�%�M[��W��]:���J���Cu�(?�M�Fm��rUF��T�[����J}[%�Q�!����y�eV|���J)��i�+ǭ�D!��U�i���NM�}̤p�����Y�����?H�\鐁�\&�"F���ɖ�X�^7!I^�C�}.�������^O�,�h���9v`=�!!. �
f�=���?� �Ck��z�L��jU>Y@ȓo�N��kJd�+��hM�V��2(1o�XΒdQ �qWmS2=p:�����}^���h�t�T�k�	��E����#�Oߘ짍>f�0�PL�>=���������E��%4�L#��#ey��(�p���9wC�J�O���NQ�.\�"������l��1���*T]&2<����\�������	 ��#W���wpm����`6�/�U��(4���O�D��䈳j�~[�nF\?[^���bfE��K����MSN�"~]�3��G����b��fk��-H�{��'t0zW���|� >�&U�∏+��pc7:z��g�ޛ��2�e�����{?ݜ?�����(���7,{kn� m;�?���������=�|y�*�:�+ �V�X��MmYEs��OO���tN%��ʹg>rCn68P��S��rӔLd�Nݞ�+�C[�y�{�xl_謗�>˿��48x�U��$)����y+���>�E����Ы�m琸V�;�J�-%�p�C[���x��%M�S����ϖCB�oK� �^Y�"�jү�dT���5�`}Ŝ��I��4�xpքu��S��-ߜ��P��j.��������@7^V#��}n	�z1��a�CR���"�`D߬�S�g�}������k"Pͱ�1*{hO8�LQ4E�EI).���h�ڳ�"#�!��B�O��&��� O/-՛����R�]O�5��a&L$�Wkhz��T�N?f̄����͗C�&���|�'\����!E8�N��n�T�V�Aaz��v4�������C؍ J��y��T���2�q9<���L��lf�Lt�U��ѓ
@c9e�<�0�O^�F�˥��9�}� �^��B�Ē=<m.A^����ÇP$��P�?�^l<��s��=s��*�]Ӂ�����n��@��fѕA#A= ���Y��V��:��X�~�����C���2�E?N�9|��0$j�3�=1;����\4���S�mE�Ľ,߷��:H��[¹�N��>xz!Yq��!���q씥;0[�������w�o��[��.���Y�Hk@�s�h#G��\��6NJׂ>���b9�Mg�?�]�,���f�x���ܦ��q����woǕ�scԁ�דrU:V�S��e:=�;*-0���o	��}kBQ\�y0�3)[8:i�,i�XlxVHYEB    fa00    1910�8�"#惦-t�d�!� t߳7-ܕ-�R�a�jٮ�R����ش�M+���^�m=��b�f)�ɖ�٠�4g�T�����a%UEx�C�������(�҃C:�/1 D,H�2�W`1c~�W,T
�N.ï25���W�x��L̥�<H&<(&�n(hl{�~հ��6m���x�e)T��Uς��.�%D�ұ��k���AG	ݐn��k����ߵ �����n/)$Z�����獬�+��j%n"�f=x?1��@��ݼY��C.�XV��2q���������W!֯�����X?:����5ح��k�r|u5�r�xM|�&��u�T\ ��h��'�\Ց�+<!#(�F'�r�����'�g[īb�{	o�u�戞Dԡk.�8�ǈ��RU��$oA�A�?J\'Av��X&ٍ�/ך��4���_�i���VpM}8	��+���Iʚ|���xB��iw��\��㪕�jk��<����Y��y1��l�#>�!��,k!A TJ��,M/�$짻/Y�W�����r���y���@-��(���.���C񠗷���ڊ�������D?:p'T�ֶ!�s���"}_�镚(�R�K�Ŀ8T��ׄY�J$g|�!~R#��5 ]�j9	l��p�0��r3��(Jⴟ�8��a�O>�m���0�Y-�px�g8�X��3�
�6�.�#?/�癃�L!H�ǌL��[z6ڣ]T?��O/kH�Sc2������P�9���7�h�]�o� �iP���{ܗ2*�֔ӿ�<�ߕ�s�"m�"��'Fy;jW��p^�� �3EH�c���*s�Yp]8@��;��hr)�2H }Z�xZ%��KJ�ϋz��o�9-	 ����Il�)�m	n�����M[.!���t��辆�\��f���m�5��c���D��51����ޘ�9 ��H�-�?X	VM����3
�J�,���h���w~Z?��/�dZ5J�my��V�fZ��x�uIEc�ݵ��p�-([�8P�6�'7��p=��Ķ�g�6ϛm�����uM�ri�$� g�=�b�\��BX�0�~���?�@Ē^�"�f�Ge�f�3��n�����Խ)�ԋ�q0�D�Sn���Q��M��8=��Ϡп���C�yO{�/a�<�f�:�"' u����������k��z [xU�]�[S�^䛳�QYU�oUg�=N�㈄lq]�r���G���p[�x,4`(�H&�M�{^�,$#���O3��ξM��8�[E� ~���@.ٟt3k��|��9K�Whrok~���	�{�B=ݯ�+�w[��\��g����Q(�$��I?�`����GC4E�N�0�V/�Y��D��{�49�qg��6�'�E��6?Ykm���UС����f)��"���M�h��O�@�*f��w3���
�6�;�f�G��&��zl^�T�	���h'R.�:1�'C$��,HÍC�7{�]�Iw���[D5���ED*���1-��@^��~	�5LS��$�qU���"p{X���X�i�(���h����l�x�9�6�ntγތqC�_a,M#��[x�8��"h$�1�t7¥���nXE�M����R�	z�FX9�0N�_���l�q VF3�,GZǚ�^�C�p�6z��#G�CfߌH��{�]g+�\���'�Sh�~�~���"��z@?1j޲���硨|����E((��|�����>W>�&���oz��k5nΖ,�'.�3�Q�vo���@]���|,w�~��}�W����r�dE���`��fݳ��w;��Hz�l��8��*[�{#��5��s���b\�< CJ�����zu���v6:t<^���*�[�Q��㜄��Te��%��b�i����]`��Lm;�����M�Ӆ{^@ L�*�ƪB�z��j���2�����3G_�m"ta��Ns�{�5l$}��A`6�(�+�.eL�Z\2F��D׵��6�p�; R�e��-^-A�} ��S�r�����P�-�����D�H�t�q�����:�wֲ؃��47��������I��Y�x��QBn@�4N��g�[}�|=`6֜-Dz	8���\�z�o�ȫTo��m������$Y�[���?ypH�;��"�ۖb�����6��:���qQ�(��k�y�٬z�U�|������R�9�k;�V��#.�aG���pzC�I1xk������3����K��B�8E�:oz42�U:�����<�c0��g�('���SL1��߃���;�dBE�&:���ih���F�i���5z�i�`w�ȕ��$�����-u���t�W���#��s^#������W/=�/���1�B=���8�P9?B�a�j�	��U�D*��k����X�s��R-=G�Mj׀�>��+��'a��_�4^�O��n0Aζ�?�iE�-6�|����zY�
��׾l��r�3\p��'��+[�����JB\D_O@�4崉�;�����C7��Ȳ�AP�VITDw;5=4�ȅ�F��ـ=5�m���I93�\�uĀ �F��ǁI�骰[���8(��g��U��ӯ��L�&2`�47�Zs9$Ej$z���q����Z���n�-*���>�h�S�1®hOH"�h/�WB�Kl�"���2��,2Mi6�5�١naP?G�Z��?ȎH@�?=��C�
:�Q�n$o��%������5���$�l���ΆAp��!A�H��J�i�zD���0�e���rN_\��nJ�Vbk!4Hˬ��ʙ$�O
���Q%�2��/qK��&&M�	�d�We�T�}2���H4��[Q���ܢ͢�o�=�u�X����y���W��cМ{43�wɧ)��"���=<>J����D�Uz��3����-�^��s�;��������
h]�f�xoo�kxгw �������Wz�\S$a�d#Z�w\�����D����� ^��U@��0�|r$��a-������?��4ߩԍfѬ��Z&�ޘ1nFjF�[7�W��a��i�/jl�/��{2�o��	Q�Ǚ�"��K�ݾ�]��Y=��ڹ^��5�T�r���Q��ȩ��_� ��QZ�	�Մ�4JF���jfޞ�C�k�Tԫ.,BoWj��p�w�,�Tn>ƴ&�r���]��T�p#c}+W�!��l�����Ε���{v>�3r��?4���L��C��E�{��_���iKm��	W���^���!&�/Tu.��&�Xp��������Qښ�W���V��nC�*�8b�L/h��I�e���af���^�~${-)�)B����)�ܧ��-N�t}xQ�?�4�#�l��߾�9�.^1x{"�k�гH?el�7q�Z��/�s;�إ`���'�4�4d��!�����=�V��x���K4r�|S%�*���b�(y]m�4��x6M�N������c����ߛ�5e��Ȕ�����&LO{^�1�u7`�Sy2bi~�����h��	��?'���^|�.]O@ 6^������C�O����f�Q�T���(:�<�I�k�2'�-��ѧ�����>�]��"Q���O��� ho�< ��^35����!r���kWv�It]fUqܶ ����o�|Н�t^�w1�t���P)��3gC�|�;T�{��c��=��t��X<��+�ߊ�'�+~�z��z��D��,|�݈������:�2�Zs�xs��o]ܔl
�>��&��2�?Q�����h��!���ow��B�����z��#�H��閒Hrn�q.�L�a�u��ܬo�=�{��Ǆ�LEH�~�S��I��4�h+�-�H�î�������4\�^D��A���Ǽ���n�@���	�kDW��>Ⴭ1�ǋ*i+��uM�<��F64��-���տ6�s8�K;a�,�����X�t0��Ce	#tc�7f�+�S���Ln&<��d<
�k�����ֶH�xe���9�r��E�����]�et��H¸�:������;l�Ge|�-�{��aFӆ��!s�_�����+ǉ�D`4M31<��ٌ���h�,���G<�	�׽�>3�I�L�Z��]�3��6!��blZ������u8��
1� ��t����J�D�����C ��;*��=Q(��f^kp����-���A#ܳR�����٨�G��X,��7'��	�2L{���m����5�D��%ByJ��Al9\d�8�L�}�͛nϤ�����Ѷ�k�~$�SA�l�����='��\���`ow���Z6|o�Y25F�x�JEr�gX�S.޴����Ԟ��s���v��ZC����?FY���e��oV�'��}��u��,�?����NH���	��p�ۑ�'��1r#��n7.�{H�����Nh�i�e��t�z������jǵ���P���b�q���=�f��s�s��o#��"�ߘf+�@+Q�ِ����W�ei��s��$T�4&"����{Eja�����ƇV��杙\�c`�3��g�d��=�E��
�pء�L�nۢ��~�ԍE\z3K�iyp�ZK�.���=�E�lyn�I�R����0�u��Pi��"����u蜮���q[%}��44���� ��X��FH�Ұ�65`K�E��Bzj���:�g�n��Ь��S����'aB�B�3BLfS4�Iʎ�lc�:_�s,�@^_���F �-�$�i�|~�B�i���,#�μ��غ���FwW�:�b�9=�{zT�+�����������3�}�,�9��9%*	�/�>����&G|Xq��o
?��H���Q��ڊޛ��MTڅ�c�M}����o��� e�P,�e���!i\_�CZzGi�,�#�G���Q
����S&ǖ��Ĉi�7;�\k��V�������Qr����eE�ȣ�i�������L��}K�Ө�wn�e�n���s���$B͟x�)SP�3x��Z�J��>�d��:�Ҡ��YcD�A��EQ�a�nD�@!U��z6�EOfK��݆��,��k�~�%�%���%��"�z,�k0�I��#��8�����S�ze):�����S��C�����V�������S$�QҶ��]��q����-I5�! ]��5)��x|={�K3��r�P�w�.?+2�ǫ��m����Pٙ�O�B.���T��ך�m�4��d Eڏk@�7G���j�ګ���fZE�=E��<
���}���Hן���j�&`�P��� �\�م9_Y
��Ib;�����
N>�䛠S�����,�nJ�$���*WL�����~2x�&~��pll�3�z}Z��
ϳ~�������F�d.�om݂vFw'���]���Z����%�TE5f��%�~�z)]�cNkr�<x��Y�o������6�I��[l���ʒ���服�'H�cY.%�{�s>u.A��b�����(K��<�<~d-[�Tئѧ�j�>��A��0�9m1�F�v̻��ܷ�����>������01��)9iqpᴇ�(r����2���z0��̓f�l�W��i7�� F��M��)lk�m�|.}v�b�)����[�&[�'k�߿%�L�������#$�O����{��1�aq����ya��u�I��ًd���au�ћ�UJ�����M� lpR�	jŐ�Vѵȇ�.^�[Z=
wӷ_'����xO���������N�0��w�;�Ec��������X�r0��a���=;�δ�&_�ܽ��l� [E�*��22!5�v|Cb�0���g,2)6e�@��U@	E�~v�2���=��.�+�Ƕ�9~_����P��
.���_��y�� Z�_&�RlR�V��C1��:����x����*�@���lT�O9=�t:�r��M��
|���d�T.�Ղ�r�`/eF�r�7�NM8��p����J���aa理+q��|�ע���j�F5�Zk�;u'#�N���۩		�̅�I ��'AZ�9��4V�͜T�u��ۙrv��ҡoƫ3��.*UB'�ηNf�5V��~E��H7�u�G�-�d����\(� +I�m��-؋��A�5	%v�xU�ƅ�.V/����yI#��3��YX�}׏�8��A��JA���Y��� xKk�ѹ�驡xW��Ul�X���Ԏ{N��WD@8��(�������8�2��8�0��A�t����>�[I��UqЮfN|����>U���fF��~_>�G������Ԉ{˽�&�XlxVHYEB    fa00    10e0Jx�/E�׭�m����i��NuuQQ�d'O��^���y8���2�z��kC���h!G�$�/a*�u�+�+���=ڋ�֋{�p��&�7Z�A�L�Ay���0�T�l�(�B޼�����2,��#�ZI�A�K�Hb窃�(��59C?\�_9i~cO�&ц��w�>�	z�YÕ�>^y*w�Ɋ�:�h2z������:G� �V�<(�+�9)������g����D� �tvBܪ�n���pc��ljz5
Yz�tм������X�h�.�i��t�����g[�/`��u��{��уx'�!�u[�t+����s^Q#4o�ؠ]�:��~��;\/�Kx�I�h&Wz0(~u�<��Xt�̧��b�E�m�J$K����-[�7-W����C�P����T�X� ��ZS�ܔ+�5�$AN;!�̪驙�ݮiZd�	}�����.��h7��z�&&�R7����.��*ҙ�u����-{�y>?؁xΥjx�l`j6]W	>8^jͥa� B_�L ���g���<�׸nVD�,���o6/q۫�� 
�8?�=$�ш��p�Db9w�F��^�O�ު}�[[~��m��l�����2~���!)N��̀A6�t-���!Ү�޺��҂�~��@����,-`�S�\��K�|��7�eR�A=�\�O �s_֮�zJ��
Q����)���#
�:`��%*����|71� P���sqߡS�6��A�
B7�ҹd���0�Ox岓S�Q�����.�r��m8�dq�n��N6y���)��������{,4�>����w�=m'�ٺ6���(�J�)��=�8������c���m0���*�W� 1�������M���q�a�|�FRԒphs�̒oe���I«,~���ִ��Ȑ6�^p	�9��R8�O��t��\8��q�(+,��	�����DXC�{L��8�󅡘)T�DE >_�:b���=�����O�ˋ�����7vEΉ���L/���HɿEA����H�'\�ۆ{�� �� 4h�nlZ���󯙌�0�8P�WCJ��\f�ݞ��@}�Ap�l�unw���o�DK�z��	� U�4tΤ�:���D�Mq���$���ܾ��8�R5įPqу?]z�Сݎ,��.VAer/��0�,��^H�Jx0[�4�1k�U�!5߭>�_�fo"� ��fV>��sOJ�yj� ����|T�_S)ǲ_���^[�+��k���@�ŷ�
��+HE��T�}1Ҫ�g!Y�<��T�8�Q&ޢ���ƑD�Cq����fk�8��r�ۖe��I~BbG�vIYkreS��:ş��z�/H�U,k���#��:�rz��$CҚ�ҿ�=-D�vç��.t�J$5���V5�*��і^&��
D��k���7=�<t"���\ՅT�,Hkq�D"�#q'��o�8���ixN�x�P��V�9�:�u��	�����Ga��^<VRu/"~�D�F���S�,�����Q�^�T��A4Bˆ�ae�� ���Ȣ� ��!x Q|hx`g������̷�x-{蔟��?:�j)�_#�IZL��߳%Ȉ�D���@������qJ�LO�#Y��!�ta�����hPؐ�R֋�f��Pg#������q
Qa�2�#h	��P#zv�?3ծ��A�F�X ;ַ�H,��x�,���D"�m��e�;�{��� �s��u��&�A*]qu�Q���O�eM�����`)�S{�+�6�<W�M�a��pT��rq�#u_�2p$j~	$����*�qrn�n���(��3@q��fB��|�����8'�΀�=���p&|%�\��襘�>)�E%�R��;qx��P�36Ѩ$�,Y��x��iU-IqG�@�k����u4;t���~BCL\�F��5��S���׹�CI+�a���el}�yM����fY���<�a?aֻ\��sL�8�#�?�!\@��ji�[diP<D;V(V?s5hnY'��%~��vYE�3����a��U�s���L���9����	�=\3<a�/��`��B��,�ބ2��Y�Gm����wf9�E��̹���@�g����SH�F,ev�$#V�_l�a��d��
�Nv0Z��X��z3=д�J=M��T��W�5M�Ll�®V|�_	V`(t�]d�/��H�K���������铋����gW�dJӌr���S�@�x*�.=�ݏw��6Hu���f��ce����w�1��D͐�邻�&OrH��(a�m��bR�;�A�����srr@����|������F?,#�|�l�)5�3�Ɔ:�ˇ+��롮���w� HX����	Ȼu]i�VU8һ���s�R��o�ן�p�Մ�^�4PhG/���x��`\k�;I�Wc*�&p:�A0�F��!Ei� K�]��<�� }�뻓4#b)���v#5�K��,����CF�����c�y���Z.�b|�IMZ	��'�.rqx�������*`o�ww]NH�w���=���$����ޟ��(ɋ��a�ľ�wl�
]6^�Ȯx�g�%$N_#�5(#��I��˸o�˓;7�PN��M�T��:�D�B�G[@/���{�kP�,��d>(f��9-{�w����:�Q�����v��F�6�d�Wn��O7��������u?g7���rr��"����̯��B��+�KFI���p�`��D�����]��-�~����_���x�㘱�_N�Ҥ�-�����(|���n�)8&��k�&1L��V� G��Z�� |��Ω��AD`�SKuu,Z_��9s�R�dB�鋄���5!&��HҩGNu��df�4��-]]�&��o}�ҙX����u�-�[��:�g�u~������#P)��z2�,��"}E]d�/ n���YS�}���(eڳ*`��H7�ktE{��Mp�\!�p�����](٘��/n
����W�'��v�Z�ATI���T�H��r3�q�D�|��z��p���i~.��ٴ�=������~n�}Y�V���ZxE��>V�����-����I
����;DG�{�n������ ��<���$?Aޠ8E�G%�[4^��I�H�.�^�jw�V!�	H����$Z�s���v�<�x �Q�m=��q9���4�7��`����`J�OWA�y�����zvų�-i��E�Ve��V8��cw2�u
}<�z<ܸm<c;�)��@;��0����!�y}�re YST�}~oY�k��r���E�*�kl��q��l����N��f�YH�r�����
R
����Z��b���b#��y;`G�o�w����fP�&�:!=� �6&T���-��Ѷ��R�|߸��#��բ1�>k��,z94h�����s.C�2���{�)"c4���q�f�5*@GiM��EU�$V������.�ě�}t�O	�������%{�Y<�Cƣ&yl&zв@DO0�j4g+�7��'�x�eP�X�8�1��
����n*p�J̒3X��eKm/���	��1�nA}^��R���7hzVEE����DÐ[As��+G�t�5@菒DI��&C�w���y���������ʖ��&��p�Ƚ��v֥GG�^+%���r&W��#G)P5c~e@i�^��n��J_ȯL�6<�;aϡ&;�匙e��s@B���q�B�'����z�"x�K9��&��kF�p�����tKd���-7��k粮�x<R�d��l�%����q��!�WB  ������G>��6I\� ����t\��\Voj��t�%��b�I�W�[v��|��E��"��{���60t��0�!�U�S��*���܉00`��o������	4����=��Ē����E�i�s��56��~^���r6T�Ih9��Ȥ�Ϫ0x�-8%�'i�	$ϋ���!ERu9�*Kk̍|�r2�l���~%c#u�y.	+�אwm_5�d�8��v#TD��$���~u�_W����f��J�k^K�3h�ý��ͨ�O�Cj��!�f����`$���G!�:u�Sѓw���(^F�d6,�+{���1��xR�GY)�e��q6�%�j� Jg�g�p_��ݰv"�聃�"�j���,́�:#t��xrn�X�&pM�`y)Ѷ�c\D�������U�Lxq��1��?4c5�{�`��S%F�]�"�XlxVHYEB    fa00    1860�9����õ���a�����2&Q�u��p�ULb���h��\���?B���`=1⡮��o�
�����vLK�����#��15�7&�{&d5�\
�ϒ��t_k�@�_�h���o��%��M���8� X���B�6�V�J�w���oL�%���дw�
L��bVW���?�k���]��/�x�at�u9�cWd�/-�?'�+y�H�ye�wB�
E�/��ç���P�\J
�t=Tt�s�W�K��J�e�	˳�^���>ѕ�Q��`�(��y�;|y{{*J��K���ܳK��h��&l��'E}`�;Fn� z�!�=i��%�V�+��/T�c5�f#�ǂ����Q�X��|jT���z!n��|�Y"��D���૝5��7P���2[
2$) �ʳ�p<�铯)wd0�?��&EK��rs�=H��{�Nb�8��v��3�42S�� �j���vB�[E�:�"E��m�8�i }��f����mǊ4�?(r ,�6�lџ�4~7���'���۝�?_�P��V�i�ĸb�t<�� ���AG�� ��uBD	�ĕ���ܗ��j��h����y��_[�Y���D�SwV�$9��:>43�Iu��U��gNj�T=�D*_5�z�����v���ճ�]�xj���!I��NwUD��6�LBH��3���L����ת��)DJ��>�|
�2��U�w�b����G�n~��B2��hs-�}<�2<0�����z�b$I�AM�2������rZIT	9�	i�6�k?L�9���]1��S�X>I���� ��h��w�S �$�,p�F�0�F�����F&��N�N²�_]g�����2���3��u��/i#̹M-���y-�� a6�}���y+Q�P1и4v�gs4G2�3��w�X?_��*��]��1�;�B���9�/0�u �H�5��V�CT�J����sׁ��)K$3�P��Uh_sPڤ�,�PP��ԇ<��{lY�ZL�7���:k��(K?�� ;r,E7� ��Ռ��x(Q�� ��zUՖ�,B-�-Nӿ �`GR�_D�Y��n6�&a�4Q�^sw�K�[���j��WԌfx�z���7�,R��D��4Xe���Y�w1X�@"��J;;�}}"�[n�{�p�;�G�?Z��W�s�ro�1�C�k�{���l?�!�3_��{�����Fh��+�T�-�v��&1��O�M���-b*}]����]�9�X+g�c91�tK]$�A|h�����ǭ������!�br�j� i�#� }�*�e����*�=C���E��5i9/�&�~P����]�*zO�N�!RC.�_י�L���GU�
���0D5f������b�!��s[+�rj���}����?a�-<�+�M�-P2o�T���-�\M�3O�O�X�Q2ԫd��Xfb�P�ia���٭Q�a9�@�6|�2�ohb���hD^��8���C�Mt�S�����!�֦�it�v잛A}�E�m�1���Y�`4�ki
8��0�������ߑ*�1��m�6�����m���a�fC�k�Y�#�G9s�R.f��S��"_]H^M�:�=�s;���u�ob����)C%��OU�1��r(ZѲ�qu`	o��'mJ=m(��#�b��������Lz@�I.�([l����[�uɻ�,�m�����n�h����S����(�I�V$��;/b=\�������8/qг��ul�Q���F�EG��h>W�'�/ؽ��
�(�t�{̅����ӌM����
� uC\���%66�Ӎ�}c���F��A���~���� ��-��"�j�~�&R�D��FU�ͨ�x�_)�1��rn��~�md�����6g�l���k�RP��FR��]Noȓ�yu}�C�(�I��?�}K��BMW��G��q`�Q�J�Ң��oo9k�<�*l��c]w�>�`jCH�Νт8g��ZD/z�]&"�Ϣ���52�2����&M6&����Rb�vO�"Hc���7���(�58($Z
�{e	�XN�&���5EgJ����MmK�:"�f@�a:wJ8���(�g��y�|F�#Km��>���S��VxC%Ns⼧��������Z�Rզ���[)���;������<��]�[V�
���s�g�6��Ɍv���՞�c�-;\��[��H�W�ܬ�m��?�&�:�p����b���F�)��k���/p��dM�9�e&x��<��.삘F7-"��QZ`�xS�shv�]��,Ia\m%�!�ׇ�����u�/�mJ-^�Me�z�:Ʋ)����) L��T#�{�M笾�2�� �8y��Ȁ��q@�b¨���z��E�yJ��0'~c7�&���	i��8���3Pc-ԗ_`�&P�'*< R�����E�f�|��Y�:�T�E@��v���* E�)�yAa/�A��=�S@QS�))�f����-����:���U_z�eft:���q�]�9�p*Y)��D(�S��ߟ���ܰp��lj��_"`x7��EzK���*W��y.E$o�?�M>.�ĎK�W�z~n�\��p��`j�U��*$��:�ˆ7ᤄ�5N�<��B_�w�6�V���"�~��J��p85�/�0�>��p_.\��}�J�ޏ�T�G�&t	zd�̸��pa{!*A�����`*z�����5�بoCN��2'V�ۇ'��0z��iE�31o��6i�?�ó�R6L�� U �q����- 8���<�B�����(>��R�b�$M���	]KX��q,J�_#3�����z�f;��
���I�?�D3������jI��dH�@4KNB~N�>�t�/C �U �~5��mq�l5 ��u�b�ͫQ��
�M?�K��J.G�q��ܤfH��B�{�~����v�f�}�;��Ռ�>�P��x�;u8���q�����8!�(aP�����.�U���ܼ�e2w}j��"�摴���zdާ8���XE�g'��]�D7�5�-�$�����>�z�;,S�;fԸ��8���kݠ�B���@�������8���K:��.��MA���1�s����,�em[�{�|�����ƒ�gL��I�Գ}��ao�M�Y��Qh'��F6�G@	{<)�D�[��Y��l:;�����͟��'���k�/��$���OҚ���-�"õ*I���=�w^�� ��7,]���Ǭ���X# ��d]�Ѫ��ȈS:L7 <��qQU,��H�x�Lx���_)_D�xw�ͩ�`�y^�^���C�{��oh�\8��{NEG+֍bV͓G�K�*�a��Z\�蜰_�h;���`��}�M`	(Rt� 9�(�gV�/#���:_��i��LN!KX�� �e"0��(v��;sӭ36������o��l���\�53~_c�NH~2NЈ ��I&. �ۚ4E��̗`�8\Nd�}&,�dT�k�o�����OG�"N%�̿��g���nA�Pl
�^�k���֋E�d��C.��wAFM�t�H���A����#�7��BtU��")m��'F��+��j���s�cMM��Rf���3T�'⹮q����I����#Q�(Z�@lO��/CPBd9�
��Ae%�j����=$��:O�	XUj99��V���{nPI�HA?GB�g��y�C����^5�i7�t�y��������o�P�eρ0<W���V{a�z��1��Ll����Q�)ܛ��I}��m������v���M���U��n����/���{��ք5�Ν��Q ��ȜsvҵIE���ؤZ���<%�a� ��Y(����N���ڂ���n�Y��Ia�Â����'<5�T�dR��gr�΄W��!! �Pxy^�@%��Yκ�VƲ����r�rq
�����@[��=K����9�
'k�w����\�ڰW�"��Б�>	#�
�oS6@˥�D?c�m���s�C��̐A�<�9�?������)>5��E@�
�^�'�UQ�A�"��LI�\!�Я*�����F�$ss���
�����,w��
4�7�'T�%̣P�L;�����1T�Χɹy����)۰OG�T6��ie1&��)C��i)	9���rf2J�B��t��K�A]]�|�������2yI
Bu��'�J�zM�`㼂W�z��'�[Ð?p�.N���<�Qܦ��#���t��N�=��KW��~~�i5�'y�}����i�2���v,�y�{�rFv�<�G��W��E��q·fR�s�ţ�zc��ؒ���������ف��͎p:�iΌ��A�Eԗ�R����B=�M56|+�� !��1g����[���l
&ymB"�4]b��Ϥ�~RX=��OQ6�k�֟މѿ%_��Ĥ3jH3�f�}z8���j�~���@�q�7���`�hc���یŉy�{R}٣x��!S�ӥ��dcB�Ŧ���V1Qs���E%s���?�a`9֕"+@r_�I�1�[�=���d�B!�2�ڭi��7�ޯp�]��:̊��T@@xC���ݩm\��>}6#cd(g���c��N��ρ�q|�;mv�"X���s�)��x�?�T\E3��ʜ�r�Wʟ�N��\"����,����<����:יMyś˽���T�FK�y~5��x3�k����t�!y�p�n��?�)I-�W	�1ǆ9=�,���GD;�*�׏<���Ѷ����̈́
Y~I�J=x��"To��!l<d����6�K"����HZ�R95���A(���čx��{�̆^���η��qW�O��S��%��7M��g�z%54��(.��B;!�67�e;׳��P���.l����c@�s&���>ֈ�w�.�'�\.�����ҝ� ]�r�����KC.�tJ�����~�l�ۉ�*��՚�v熾1k�����z��t�0�����ֲY��|C����K%E&�8��;����e�Ħ�ft	d̋����#mjB�tR��J�'1��O�]yl�"� "�!F�	��K<d��}o����&����������,:%�h����0uf�g��r����މG�:E�|�N&�ϖ��}��"p�����Wծ�A/�`���cڤ/.��z��L��z�c����
���|4h��^��#[i9F|U�g��ƀ�h#����s4�4]��J���ZY|��Oa���_4	�(�>3V��� S'�8k��ƻ%��s���F@��Dv���p3-Jqw�+ ���(=z��������������x��pz�Z�W���~"�4�	G[iv��}���=Y��&��Q7�3caN�~���Q��g^0N�)@�ބ���鍕L���ӓ�q>m��Q����j�zfM�+�g�F�.�|���}:, 4X������"���K��r|�)o��y�kX��5©X|������H�0~!�Cwz�TOg@[��΃"��995���x��l�!ek���s-�H���}���0��y�^KS����]�$q����G���%u���v����"���sp�ܟ�������1Ef���e�<GT
;S�$����vdB�d�<�"S_a'�y��z`8��c��y��� ���DJP��PW1�S��5<
L}<Y�;�>N�S��@O�a�>�S5��ڒ50�3w�(�L��I�R����?�vh��������}�]z�^&a�;�w�E�#
�{����n`�v��c�FC�gl�$�������&��Ej���4ד�oh׃��{�q)$�K��Q�y	Ok��j�!��K+]�A��5���4��-C�z��T3*FVR��J�����ج,�* xV5j�����_Q e��y����^h����a��[����Y�^��bay��L�Yʘ�35(\�E
��w�/��4�P vz�p�֕G�"^&c���M�mʼy�����\1^6��x�0;�K�Lh��R�Ӯ=<���<{������H����G�@�����r������!�b�[}d�Sq�pc~�R�aw1�S� /���"�P0�P�.\r�����*�`.�k�ld�B~��<XlxVHYEB    fa00    1720u7����v�k�UtEI���w2���t��w�v+?���f# �Y-Ϻi��B�͆�EW�nE����|���f�[E���A]w~s���ޠ���2%�^����������B4��[�:�����ɷ����?���zm����V��(svE��9�C����<�A�m	ؗ\�v�p뫴����[�@�י���̆�9��@rn��R��q#�g��[ڐ����^��A�]����@��d+>$#S㷺�0�ug*�00�cF_���O'�@s*k$�+�yF�c/��1�%Y��	�wd�r4|0��>6&�C��sˤ�-�EL�'�"+��.3G;�/�N�*�o��<�jNS٭���Gy��"��_;�ʎ���y�E�.���'jow��X�� �s��"mj(�{��w�d���.c��@*�I�,�V|n��q���P��DWv*4f�r����L�@I/�ߔ��1<��R�CSw�������H�\/V++�+�V|���sH�q.���J?�o'���e+�G�9�Q�˻��`-��KԖ�)z�f��Q��XC�x�
9d=h��c��T:K$���f:ih�
�Q�D���d�'�<)U&�x]�T���3�8R��������.�7������h�shEDaB�'��`�؟������Ҩ1���'{K��&tF��xe�QL6�+�����#]	�����n������n����P������x�O�5��З[��_��|�Y��Ƞ��8hJ���_��Zcڔ���Y6i۟�=&K4Ľ�q��Pz�M��4O �i{ mo.T|�T� �Y���D�w0v���&I!�z[v*�\��}uso{��C��b�L��G�\��	D��4@��1䐛��\_����Ij���	
cO]V(����>C���뚿��!P��x�U�߅q��A�;mS� �^{#����AC:t�b�!�ʤ+�W2=W]f�]>�#U�Z�Z�qzZi�ve+BI�=��I���e`�R0�[���|���߹�3�}���ic5����M����\�_�A���Ժ�!$���F��%yD��X��dRC�N��R�ve�`Ww8��y'�_�	1�κ(�98e�� {�~y�b�xz ']��Fy�& ��J7��(��O������be]�ۭ��-��]m!�h�	}T�����~߄0��g�>,~^�7�Ȓ]跲��Fn��4 b�:�l��l�Kd
�<n�N��*0�B���������%n��xR�BQƓ�L��{�~b(	6�7?��3�����~� JA߰�fvC��\KC�U��C���⁆FA#�O?�<%����װ�cΟ���YǺFQ����	R���P��a"�W�#��������xo <�bth��A�L��"��Ａ2~��VjR��:��|�K��{c!X��f��5e	!e�tބ'1freb�� �p}LQӓ��<�� l+/����n� `�;�#8�F�ߞeB?$���1%���"��6C��4u��0���Ü���g���5�;�m�Q+�����8~�M��#�w݈�oDP�a�X��o��N\�����WK;��x
��̂>��<o� ��3��raIA�^���NnА獑щ;@L��}g��#N��_j%4�<��,�OA�PEKd(���ь~�A��a�r������!Ƽ��������@��x�����Z��@�� �8�E��Pn�?����6��!�օ�0��%���
X���N�=_����g�ƃ�E�
m�_^$��\~�w9{�U8`�RzF��6\H`�.���>��rk���Og�⫮���q�LȰ��N6os&�OPL��7y���P� �!�>xV��_��BS� }������-�tr���K�|�Ԭ�ʈi�|��mȏw�k1�ᏀJZ�8��Վ�$-���~�7�#-��JذI3��z/Fu-���ĥTq���"��Ҁ�����f��G}�o
%�B���j�Z~k��_>\��ޛ.�܋7��4w��5 0(��<؃�������X[���w$1�a,�D1��ӓ��8�
%�������h8���L������#����ZWf3�v>it7γ��V��d�P�Y���0"O������d�ΧH 0�y|�|q�������)�ݩhˬN�4<��,�l��($�n��	�P3T�&�}�սf�"v��\IT�ޢ���-�MA7�3��_��*��r�%�]!�r�ߞl�E�l�!8^G?��S*���@�s���y!U��=W�Q�+�z)DJ�/�e���`��ú8xB�I���X�XiB�k�\�|�C�i�Zt܏�#hH[�%�����{�'<>��־@.��Xbuq���;׉|�yr�s��.���&�]
:Z�sQ�Q�3�y��k��3*����5T��|����?;�T�?����G𾗤g}�G�B�=L5&,\"4]4�Z�e�^|�/ P�Ӂ����OH�"�MY���r�f�%�#�J�sjew t�� x��g�?����;䀧?�ӊ����#�{��sy�6���dOi�>��[?�/d����+�RЌ�Q���[��v�L��>�^Zƅ�Mt��ud����/�ͤ_���%���e��'�d�9P��yǷ-�*\�6s`�����Q���a�*Ѵ[��T�A�P�c]�1H{�w�X��=���B�~?��G��U���'���Nh��4��(��-ݬ���w-�)�#������b.l�V��i��uz��zX�,2��Ϲ�Tu�����#�D��Z�uO��vo����m3��8���hu �60���Q-!CU��'���i�t���FL|.�"�}� M���Z��O�?�����ş�28Z�@�W��6��j��d���_����4~�gOj���p�ء�_�	�^cJ��5N����T�$�鯸е��L��F�/t�xX7:x�N ��j�5}r�k���e5buȿ�q��B��#.眒Zծ��k�6�rs�>��mX�7�8�1�F	}�+���!�.b���S��g��SZ���8��S2�JI���3���@��"r�e�,�xA} ���Nb��� ǝ�u���0��n�L�$���#�O_���#m����_���\�!�)�>^���7W�������;��*�;�z׌���'�T��fw�c���pq��|D%�������3SQ�>.�v�6<y�a��B'�����n��Rڪ�`s\�Dޜ�;ow ����F?��'H�����,��?D�����KYq&�^���{�w影�?3��Tn��d(H�Z3?��A�.(�3��zj�4a�.st�ї�C{���Y[��˲&_�!>��a����1�4�����N�^�6$%6�˟������Vt��=��Gi*���X�M`�_�_	-L(�AMG<XY�����$6_d���m��b��f�e����V��?K�&薨�ݡ���i�O:��|���b�W�M×��gMkP�\��a���jқ��b�Dh
���b���QOw�{�����R��ǈ`�)|��]��M6'Y���^,�q��c�I�:4�qYM��W��[^�7��j��?RkЖ�G-·;���С�o�����=
I"�!8���{6�a�f�%[ӷ8>/N��4p
�؟�I�z���n��'�W>�l/A��Mp��6t�'��x�Z����5�g�t�TDB�1����3@�F��sS�M��s�.bBod��6�Mckpt}����h1�c1�&�2ioB� &�?��F�����I�8��Z��g�0�v\��P�l�������	&
*����J�o���f�֠�,�v�M�ڸ��*u�Ym����\-'3���q�|�B��@��|���qVk�����qxR	ۧW@i���Y��"t��W�5��@@KeJ���l����Q\�T��� ��h��͌}gΙ@�(6�a,���7�?XB��܁�_*-�nb���n����:,�d��Ɖv;���l�0b=B��Hӫ�Br��ޒW(`1�,q�T_�W`3��v������y�˹f}�<����JQ%ʠ�@+RT+�a�O���iq>e�]2ʱ����l��x��	W��D3|/��E��N����Ź}��f��*֍�o��qdE�<�s�m�Ps�ԗ�}Q�A;+��S�Ma��>�d	��Hn�9���Azx~�֓bӣxg�ቨl���ԃWB
�E/��3Q������u�XCN���E��N/��%���-��Dg���ʷ������_�t��1�WIZ?�����3��t��x-T����i��B)%SEdk�jx<Zns(��.SH�'�v��N1�tm���B�
�4HNfC����>��B������q&�� m�)��aju3���\��oT�<�+y��֒���L��$���Me5h7�8ly-@����W+�٘��:�,De�T��#L�C!	$�@����z
6�/&��Ý��&�ŉ�y� ��O$��a�{�۽`v?��4��j�Up��� �(:5�Y���<�����g
5��7{`�-���Zu�B8$|�m�F�Иi	��I#�˶r�q���e=�h�#N��Fa J��D�:���^��=�*z����	Ћ�!iB/?J$w���D�K���0��q�+�h̭�'���ŐmA���_�	�/��K���rM�L�^�����n�10�� ��T�0���gM�Yq��,��̽i�o9���&�M��
\�QR"�J��.�h�Ӧ<P��ff�G���|�7�2�
JpXc�n�>l���Z�,<�1�:�*s���d˂	δ5�1�>[���>(7:�ȯ=�l۸������t�U���&������?��((̨�7/vxî�t�(�r�Ȧj��ʙ���!ۄNK�[D�w�,ğrp�P�ic/���yn)~��oD���.�!VSaG��D��8>�qwO4���+�q�;�o�%1�`�:�~A�߿zc��ܟz�ml�W��	�<$۹��:'�X�UIJ�x~n>rH�g�	���5�`5�w�߰��M���	����̾���q� ��a6�LK~⏝:W�1��o�(#s@$��~�?K�\>$EO���u5B(����!��R��	�KV�������g*�L|[�Hi�E�L�`���)l�Nc��s%*z2G檴=Mf�峋E[��E+�~0���_�G�!���ђ\)�N�^x�<i�.��)�������wɹ�I�t��+��֌��i�L��sX`:�?�t^�!��R0d��Ƒ�:�Ä��+~qG���:o�R�'L/lXvB ��|��`�ٙ��o4[���!*%�C!5�eݞ�pO��p�_6J'��e�S:�.+<�(M>�v;��Ӫ�.�<{�x��*�"8am�����W$�I�Ip�%.xn�,	|0L��0d�S��)l��璼ٰjˣ|�K��6�Ո���}�-RC���
kG�:��^���>n��ak���@��h{��M���>��]m�Ȣ�!�t$_��Nw�.$�l���X��s�
ʛ��y�Ƿ7���8�K�����
o����aծ�O�ݵ<�|(���0�-
ܼc6�KJP;��g�i�?������ r�=M��T�!e���^�DQ	�v�~���c׶(�k��a�rJ��Lּ�����Û�I`�1����\�<+��u���(X�y�tU�y0�>U��Ew�����&4���M˒��nk^�K`�O�_-�R}�!���p�\�!�G|���1��x��U$Dգ���,������L?��k.C�	o0��Ҫy��Y�Q����5.��2���XlxVHYEB    fa00    1500?�a�vL�}K#Ҥ�ɲ��[x��I�Q!���]Z���.s�F�\h8���x0���l�O�S���#��TK�a�V�]�w�L����c,�6���y9�=-A�ˍ��!����ή4ˆp����q�đ�$J�c<��6��#.��$������-9�? �=�q��u-��}�&: l�{�.I�C��3���x{(��j�ȿ�� ]���.0 �0ޯ�����
^��j�;�g�����Z�ܓ�@$^[U$p@��?�fsKB����1f�}`ܚ�?�.=�;��#w���8�<}¾MM���9�����`��d��)ٚ���Z\T���ٕ9� �ӳ"A�+�.�-Ka�/�U�O����Hr���o�$��hu���ɖC]!]=��6+����7�W�k��)ڠ4H�šߛ�<�K(3��(=��26���+i��"%�h	Xo8Q��� ފ{��ê���[iؤ�=��t�en�� ���Q���آY��j��S���z	���?��C�λ���wU#cN(�w?�J����&��b�q>̃�1�SC��H��ۨ���9��L%ͅ����s��L6�á��l9�AE�y�Q�V��#���1�*Z�bP:�B�.��$a��Y�ZO�z���bHƇz���u�S(t��ǈ��D�@�V����H(ZU��ζ�q�`=����&�\��]a�h핟~BUTa�IJ;�UH��� V!��.�Z�uA.��WJ0�`:�#�t�[}q�_�%R��R�hVg�G��/���#`r6ʒ�U��=��V� I��װh���l�o�7I��^�"N1j벯�����l����M,KI�P�Mǒ9v�Č4Eob�>2����J���/�SN��@ȧ�����<�M�4!R�>�/����H�ŅIs���^�!�Ħ1\A���n�\+�󐳃C=8��H�8s�S��b��.x0iw�����з���W�pJ�S���'��	�PW�F+��.��"��r�U��0�1�b�
̣5�����#�r~5��|��qu�A�*`=3XM����;z1��t��JN�B���iwFQ3{C���<ڶZ�
��W�JPK�{r,qr�Ml����2��`�~3sA�{��Z�� �1��R�z.m@mc�u[�ُ��*��|ƛ-�h3%u֏��/J���8l��'�`P�Gh/+�l4?��I��h�ȽnD*F��>Ủ�D��6�G�2va��[�	�cKFjږݢ��i�$�Y��HDχ��~~���x�}�v�>f�a� �J����Yj}�2�e*��]P���8���ܩ�Ά�<����5�
�!��0�>]@�N�)�l��
��Y�s=����\(DF����kT��>��,�����M��fr%��X0�	o��N�<`��kK�k����� n��q��^Ѽ ���fY6�O9��n�U����p�	qJ:lŏ (���c.���"W�J���H�N�x_�9����].���Ȏ�
�s$L?�G^ ��1y��M�|�-�v=�>�G�?�X��%f
�G=<\��v,8���}`lK�����o)�#��ri�Q듣�X�]7�OW���^6�~Ƶ�X��)
�i�����	��VA����:�=@�H���A�v��=C�s�`E�J���`���fi���b�:b6&���EBNJ��`R[��Dk�D�,�glIOT�P�k�QzZ�!8�������me�U��(+��+�$m��lW)!��Y�������c��I�P�$�q*�t������g�t��-B�(�8�gE ��2�歁��������8���e�5'�O�y�Q»F�$�H+R���]�C]���y���^f��G��[�MY"{�!�����h��k��") ����ߛ=xQX�`k4�d7G�:K�|D���T�j���b1+<�s���׺��
.��o?3�����h�����c�����)��恮o�o,G<2b+����G�<\�v��� 5~��@R����Er�2��0|>;�%F�RTś1�c7�ئ���A+�)PR���*�W��,��Z��)���͉�vA@�R����$�KϽ��������Ub��^£o�Z���)-N�Re$;�E它k�}��y]�o�2�C:`����\sDR�n�ox=�T��ބp�D+�Ҫ������b8��~To.���O�JN}��3 Z諍���n�1�L�en�5���S�~y�AR/��?3�~+��%��S ��t��vRy�~"}Ś��'4�F��#Y��������c���2����j�?�۟ӂ��_rW�=�D�A���/����,�A���4��O��p_~0V:�zR�29��y�$!�)����P��]#N�i�r,�l)WG�5���ʹu5��?��k�����������Ր�{��*�p��Pf�{�t��0)�@[��䨿�R�b���B��ܙ���L�=rR%~����!�����Ç����nA�s(d|�ͭ�r��+0쑣���$(~I#4f�[[��z����`���grr�}���:r�@S�D��"*|�y8 �\rK&z`2
�t�.�'{)|�#�M�(����!��BA��zڝ�|�dUv?Uz��K�n���ʑ���?p�8��)�'W��h0�#��Q�tQ��xv��Q�:�־:*�B�C
%��(˞�(Ql�+��i��u|ؤ\\��
��P�=���C�#����Je��bh��:��@�`����$eT�TE'%�&�Y�~=
�-�
��ժ��S��� ��=�Hg3�%	
�7�15h��}���!�{R��5����x�2.��qǠ�m�$4���9�=^�r�����)	��'[�;��0f���Q@�xc�(FDV>kĠ����^K1�U꘳*�
`b�	�1�̤���@-,���Ԙ�^�"]x��c@KJ~*���H֋�JI$�	VB��M�|�ת��ϣUi������<��v�?�p�a;[�<��s��!�͊��@�b܅���̡/� D�#�� tɰ2[��e)��q�{������pIu�r~V�S�����J�-���u_�<�a���t�{_���|�fO����Lx��}#��z��7#����HX�R;	��憒�����3�@#��)M��S�ͪ 7����.����[��H��^�j0��7D�m��nFS����|�7�XLY��;�s����⭉�l��̆��o}ώ��� E�03�z.��KV�̃Er�և�J�J�\��!�Ԩ�(8�"��/�.�bS5Q��Yb�&�uX��i2����gU�t�4��՜��i�Wc�H����i�$>\{���璊���z֥����(�B��=���{Yu$,/�C'>d+y@ä��V�:z�㩗\Ab��Z)���\�u�j�l�Ⱥ��Tc����M��'�91�����T��;���>͜16�Ʋ�ա�B'F�E���xg��Zf��I���ӟ3�4@�ud�h0���Z����f�o��ԓl��s0��g7yH�Dxh�p���.m�ڰ���J���)74n��g��H�Y����.�
�R�.QA�V�S��������%~#���p��z�l�}��� �sF�-z�Wu3c��X�m]vV�gM���¶��X�'�,6KX��W�K�,�����h�߉��0-��Vᄜ�Q��(���ݼ1�:ª�qHG�����s��� K�+���^j���ڙ�v:����댞Q���o�B��|��sc��%E�k�ͣ����C��y��Q2HR�c�iI�ӢJc3����_]��)��(j�^��`�e��>���J9��[�<�_��Ft����.vIB���\�&8���A��޲�)����`�& 9��+���J\���z.���a�.�3_��π���ko����5���� 7���c%�҆L%WE�P3f��i b�B�k�7aOG�"�k ��R�Ɏ��r���X��G��M+��O�:�jr�Ə|�>:�8�cY���O�� Z� t�)��b��}���<7Xf�V��ُ�p{:�~0��0�0@��oW����)�v3*�����if����=Z��d�5��X�D����"v逛;M�=E-M�P������
��{k
����Ő�	sf��y��W�|�LO��900ԑ�ىTľ� ���b̀BRN�c�Ȱ�XFe��ŧ�Pw�z�-�>��	�.��|�Z_u��w-�h4��dlM�
����-��5���\7Н������|H��6׃_�j����@@��T?D���@D�9n-��Rp��Mw�R{.�i8+�9���5��$�O�,H_1�\C/�w����m�σ-��R�ca�<r��hx�c?��MMv��wWp���H�d��y0 'xu��PS_|p]i�p��;��k�^�6s�[ͼ���	���rH�i��"ʡ)I+���õ�m�yP,2)�Ĵ&���:  b�{�2Zr�Sq9�i{��g��hY&k�����,�V�s�d!.�>ȇގ+lJz��z
/;�&�>�ڴt�[\3��G-��N5��{�y�P���go���Z�U��>��j;~�ֈ�E�;:F� ��5l �V�؃ǻ�?�u���j�1]�|F�Ϙ�t|� ��ߴ����֬ϸ�mQ��s-뽓JP�}���'��xF�֚�G=���&u��ր���I���[P�P0�
��?U�薞����^�:��bʿ%�5��kq���D�M��"�s�ҝD,'�ܐ�X�����UU��?N܁�H��;�a��M莋�QM�j�cwf��I��P�f'd_����b�����;���jno�f]
����l�֞ð�\�gP�<A��,��N\y����/��:}�{���6��c��#�%�1��%�s7���H�j��N�7w?HF�<oa�_��dԤ�&P�����2"WD��S��h�i�֩!�|b9%��Ҿ��a�7�q��b��\�Dﶔ�9���,��p+��p�������s�iT����X���s�[RI�����s�ȑ�	��O�r�T?HYr4�A�CO:�2B�(BX-*�+ڭ�i ��LxNN�Q�$����:ձț_�q
Jh^�-�e"�sMÜu��]�.x _���Z���U����8B��t� �j�LI���7Ȳ���C�J�Z�I�2ޥ3�-3`���t�R�� �j���ck/b�0H�E���8A���"e� K��ۛ	��k���D,��c�,�?�bXlxVHYEB    fa00    16c0�-�f�`3���LE���Q_�ի�%]���3��Z�Z[�j}y��i�����*8�s8�5Tzw*��� |���"wò�:��o{܅&���}=�z�x�z��
D�~O�nXF���ń�=Z�Uwր�ϫ��>B�aX��[s�ロ6���!�@��yq�o6BUv�iT��+SLz&�������˫W6��	�%=�c%n#zm��ٴt��L7_�>�r���&�,���j:�f/"�+�-����}h �8����#��5.e�:x�:�	��B��<�g=���AzJ�#	�i��w~*l�\�T̫Y%��!�R�r��XT7%�&L�f b�6�7�W��r��yk9d̎J40��t=�l.��S�֧C�"�c,�5鸷�MI)Y���=��(h���V���pבd�0l�I+�?9 ��$�����M�|�$�Q�����S��K�w�'��1�RrTR�c�+�J��[��5�s�A[(����~؄��Ī��8~~F?�'ݺc����VT��O��[�mKd�1t��d�.&�W�*��7 0���\���`-ه��R����IuS�CԴQރ��+��&�/�h��΄�L�Ք����w��'�n�M�yt��<�)�������� u(�&gG�N�R�!a55�>�t�d=��R� �j�q��1H�k0$E������/ ���^�xxރ��!�`���@���l0r(��'���T��e�dw�@~8�Yi��HE������0��	�ٹb��5?~8St��%9�*�W�R�|D��_�w.��Zg�~�`����U�K(<d��N5�bO��Klz�m������íN�R b����`�~�t��q+O���+�{r��+����U����$�����n�wЌ��i�\ڽ��$Ձ��Ϭ��C������i�I\$��gI����������A	����3 �K�2�}��,����r�\AL
4���'E���O��.rN��,KY�X,x���Z�tӳN����QŅ�yĺ�e�!Uȯ���g�%�&��@�3J�0`���ä�H��u\3;�F���fv�W��1�Λ#�xX�sb����ĝ-m����;���>���hun��SFNz%��c���֪=�a�i�`*�Z,c#�Q�
׼,�=0�x�.x	���Za�|����F���6-wt��Ł��V-\`�/���|ԟi�AˎG�
��J�j������e
��7����=y&�;��8l0�;FaZ,=�����>||i@D�͚��q��ө�u���Q%��aT�M���ޅy-L0j��W�P]���B�
�pÓ�5]��$�?���"�XR��CI&���G����8�����k8�� ���׀ȃ��)�O��#�\i��U���B�����Q�+�ҧ葆q߅zQ�z�i��f�en��d[;� �fHhX�i��[���P��2{�:e^��D[}�v�h�z�-H/�F��å���-��.�K�*������G_ʴ�w���-�fCw���������{���!�k�̎<��'V�������Hhk-f7�՘��Z��:?t�e����%�V����F-k�
�m���D�3�F�-{��9�BƏ��%琗_~c(���d�M��Cp�=�h����3������/�9��um��e����]�L`��$���N	�i�fK����+9��`��w��P����.���Mh���$�: g�v�G�*�D�>oD��*k�������{��1����������u����T��������Q��G���+��zҾk��`.�����H��n{�!|5�IhK# M� kS�ǚrM�$��V�8ٗS2��75���.�*d�<��Q�B$ѣW癲�,h[�O����Hg[��K4`j��@L�z`�m<c�c���Xj��lE(��2�u���R���l���z�
2�~�Ұ3��aFݧ��| ~Ǝo~P�Qh��%x��K\���)�ET	�/b�*@�KeU���Jk1�f�jb�kh-U��k��tg=�k�zTKG��D��O�yp��n�b}����=�������b��H�1e�����yP* ��^���3�s�3���Bz�ڕ4���uue� �F��Q-ك��Z
Չh��<G�j�e�eF@��R�2�^�y���0*[� ˵@S�� �J�P�����e�`�g����p٫���.�N��0N|��pҾ(�?�X���S�etLF.ô��;������K��R���I���w�&�YT���^n��ƴ���熄�<f�qk.Ԇn��h�>`��ג�s	v�
����%[y�BP�F4h��X�.ŻK��~{�����P��=l�+j�<�%������>�\ڛ��#;W2���ɿ"�����v%xO�_J���vBQ�zN�Q������M'd��`zy�KU_��%��P��[���i�E6���'��;e����3u�]	��� ʧ�wZ�P�爳QۑH���L8nu����i>���P
W�SP�6V���@�J�
QA�������ZZ-� B�v0���WOE��P��!�m��1�R��ҏH����ᕹ�:�w��y��T�����C� ��v��@Xai�b	vpBJ�	/�(�/ed���@� �����[�\G����[T���f�@?�󎕤'�ٷ��)UF�����z��>���J�ܲ���Xo�.LN�x@ɚ��0՟ SG:w��q2�V�rb��^���7)��4��E�H�#�<`�;�%W�zW�~gf	tL� j��\�1��!#�3��=�����zx[u���.\OM�bfN:˝{�$\#3}�C-��ڊ��$Ren�\�m��ͬ$��~ڀ�;(�a����*/�]������ûڢ��E��W?�H�ͅ3���bY�d�߀l2 ^����02JW�~*s���B�}�8��l�K�Q��_��GT��Tl��/�iP��9�_t�/��K��gF�Q���'H=dp2�UA��a{W�ز����}�r��C(�c�FEa�ˈnJêE.����8q��I���|���i�<�X���=S����$WF�$���n*;�"������~�ɴ7�h��TV7p���l�9Xs|XMjK���Q���[� ����o}Y�R��~�d�e����@C�����JR�4�p�%�3Sc���tng��p�̵��g��mƼ�MS��\{nW ��ࡄxm�V<ޖO�§���s̘鰥s<�A���c��۱�N�f�)d�|���t,��`>%4�K9v�M5�`��,6�ziQ�
T���D�c�ݜ�(�/�C?� ��A��U;����yk���+��C;��@0d�3�UX�:zL�7���Dɕj�rӉ�c�����n��AF L�R����RW6rղ�����
��t4�U$'���[HW�!^�{���8����#v�fcE3�x����
	��k�,k5�� 3�<|�l[�MU�&^���/$��X�>��ȃ�}��Ҋ�z���\�A�N��NT�g�z4�+f�^۟�W�[��I6�`����b�Z��W��9~{���8��`~�1�v��!�v�����I+`�(rcҰ�{�V�<\Y(���g�<�����^��}�������`���2��5(�zgEE�$�2����>[e�C4���N��]~H�m����y��j�cH���h�ܳ�V��u0pl�Bf3��X#����S�!�?��@�)���� ����g؅�cO�^&V�&%�6#]��-�u����xP��+�>|���߸3B��u� ��2�����Ɍ.|����q5$u�vuq�",h�lpU�pʷ�o�p�D݄�5�?$4���X.�p 9�|��zK�t ����}+;�H⌻To	q8�j=O�oAIؚ��e�:�L���;��i� �8���Y&O�dO�й. �ݽ՘�V �0#�#��LOة���5����J�v3��&J�9{�;+�y�~kr<{�7�8;~�	}��0����<-�f��c��̪��\V�\Ó��.W<�P�ٲ%�O����n@6�}.h:� 5����s1q��8i����Udœ+��S^5˕��6�B�"l<��Dy� ��B��x}�q�lj�a�����F�I�І�f�*H��\Y��-}��V�ʻGS0J����5y�ک����"�����w�>�-���WtQ���76G��<��0��Ǝdr�Q�ڲ�z�b���H@���;4�����^��ܗ�~���0�Ⱦ�w+��:B�f_�&�	F|T�]0��fz���a}B�'�qəd�,�R���^��b�K�,
�/ѹ ��-NɔmQ,� ���כ'!)BB�u�S���?���n7}pPB�f��~�t�g$t�	������7j�&1Pc�e����C�2��t��*�W�r�5�^$�;t��	DaY�t��*u�Ǆo�[���Ά����ϩt�!z���7�5����C�<��E���v�Jp������	��_g�gMw�� Ŗ3ӂqw��f�v�=*Q�:4�S*���{n��sV��t[8�~�r	��E��e�&oR��d�(�;\�Ƅ�;����a�uD�	�A+E���B)]A`��95C�d �eT�YTz�6�7i�ꢅVF��o�;K�'������$JNe�H,	<��\M��	��d��=x��qf�Z�삽�P���Ci��>	(�T��N�V����(�G��T(�ҽ�'�~��w�K�J�a|˶���*�����~\�`|v��(>)��B`��c1(���!MH���2����9*�%�}mM�TH����+��z�I�dk�L0;q{̉R�Q�`�Go�m?��9��o�'���f��:�~�jA��Ҟ�&P��+f 7��E���w�;*2X#�/wx����$����!���8�xHAiO�� ��{"��C�0B.�݄v������hȎ*�b�X�a:�3��}�)[����0X|gq�X�%L���i�r����p-%�`%�`�#_m��ݽM�O�ifl��n��%�������ʕ��{|,�ȱ�XX�ڎ��g���_�hX�X��`�3s�[�C��Z���M׀��{"��@����e��;}��T�},q�ʤ�튟���%�7(�`���=ݺ F���&��/)��ZԽ�B��Q�*Dy��uF��EI�/"Xp�*&�S����(��N���B��k��^�,Q%�B@PRl�o�	dh�:*��Eb��9b�c��$�w�+�6���A�[l(<flp$�*t���َZ�]�YswN?Q��ϓ	�y�a�_�Kt]����1l��-'��)�������3�sk�ݪzV�RwXZ�$y�.�AG;��@ĳ�jL)��v_2��ʶ_N��9虵ԑ������ñ��~�6���w�gŷ@�(�r澱�+]�]�\vs�����XjKb��Dhq.���y��yK �D��x�KĎ$���+� q�����G�|� .U��O8z����#����������=��X{��8�\��4��K�^�s��ͬ�+�w:4�/-�o���=C�l��E"ů�����a*�Z
;�}���|�x����δ~�Mc�BIϮ�N|���FYu��C){xy/	{��ω�n�4g ���u�����O�þ�[�-�I��d)J��v#UXlxVHYEB    fa00    1740*X͗+l��L���� #(YW2�E�!q���գ�c�ɣ���୐�s>s�>�#54JJD��t�Z�~�䲌�$�'Ɍ�F5�|7	�.-�e�|�0p^�<dM�z�q�Ō�PЅ�^�0㏿t\S�˙bf`lcq��l��.�}-��ī��X��,L��,�|����V[�=�7܅z�~�I�u��V����m;]�=F$�_1>IuK_�NKh��||=Im<6�q����
8Ex ��L�*���V'��ŭ�|��jS��"�bw)��(���-�p��շKYm�0;��I2&��}�U�	�_�H�XE��JY76E���c����I�@� �V��Ԡ��L�a?�K�Sџga>RN�D%\7��ˋ�p,T���f��L_K�SÌ�y���r����+x��%����.�h6~4$x*�C�R�kX0�ΝJ)�K,�����ퟎ�a-"��3T-���2���#��qq�����?�HM��� &�A����tvZ��e��)�ISz!�G�n�e��k�O�'�#����j	����P����� �=3&��m/o�q=ۚ�f{)������b�B����7>�IEȵs�\�ɘ��$˿FjJA�����8A�9[�]~{Ү�kPӀ���dy�������!��ޑ|���t�SF� ������65�~iLo�ܤ�^V��b������w��(r�٧�X�A�oɃm(��NMg��l�z4,�UP&�eoU&bn��O��;$��0*���'�e��1����Q����q����K�0�%'��KУ�`n.(fUź-}A���$��֍�P�P��ʑ�q��1�����gݦ*���<ŭ�ߝ�4����h��/�Ѓ!4����}�:Y�]�f6�U�?O�.S�2�ml#�!G�_�{.e��k��V�K��_6��t��&A��+a�s�"����)�\�z��ɤ��@�΂�s���ͼg<�{�7{�r��)7sy�Y�!u���NTi;���]��#B��6�t�|VbR��x�o��/�.����@�S�X�{���w^o���|��C�H�察#i�C�Z���_��B��va������u5��1z�Ȱ��uV΁q9u�B!���N��\���q�0,8�b��ڦ"&�)yN"�9p��ؙV��k�V��Eș���B����̭ʟw/�@�	sO�%{4�Q�.Va��J�@���.1��gى�C' �����nQ9��!�[Fj܌��aT��hm��TCL	0q�O++�̸��)��[H0U��l֔9}��
�-6�@ӓB?�j�.�S &�hk������R�v���Lg����#^'F�'|~����!���O>��?��B܈��J-��ڢ1tqF�'+�G��u�W`=���ǹ�ܶ��"��*!��2��Y�OԽ�b���u�[�8)mX�%)H���f�t����X��gܖ��g�X�4�Gd�]1�;��Vשj@ �2��	P%fАx�_�����r
�xHPМY�}f��bXRq?�m���|J;�����:oZ����y�P�d��oF�(��̥��7d)P8�C�|2e�6݊[��p�2��;��I��d3��A��7UH�cD<if�����Լ9�?J�\�ɭ���tr���J��fM�
��t[l�7��E4i�o���X,[Hϙ(?��y&I��J*�l�V�o����"~s�5��qGʰ���q��Y����	H�I��>�����I�K�k|�����z����,�(ie�3����U# SW���j�Icm:A��6��0F�FC[�v}�jwF ��g�5w2_q|ρ\���{�������C-:P�}HZ��~�V'8#�
���k?`�)���T'qipP�\m�*�Rf��F�.H :���6�?�gK��K?c��{kg��x���T?>�r�P��IQn1�%*���_�%�A�/��JU��흧��sl�1�ώ��;��߅��h�t��#�d�m#����!:���-���ǟ*O�5�8d��6vó���e^R��v��T�ˉ�+D��3������*�A�
3�e���@���А_v�-��G����Ҙ4��P��^�RL�
?�2����T�7�(�޶nL̃��{+�)̄�{��ɍd�g�f��њ]��hxn���'J���-L-F̆�D�h����;yi�H��$M�������)s5`5�|����JG�ω��
n�	[�e��~8�*�j�J^ ;��k;�.���ƀ�5b��D-�_���Z���$�W��.c��������-��~���H�����>�vs�=��G�:p�[#_�¯��TOh���\�w��O���vp]s�܊i�����������LS�dŋM?P�'w�J�B�9��[/�*=aIL�@��>Q� tc"N�@	=d
5t�Px��k��4���ғ�|�w����Lūg���,t_���{3��oc�WZ�JQ�Q������Oh����	��biV�}��m�$Oʪ�V'󒺖Ƿu�{��Z�΃*@�E[��nu"�AGnh{��^iK�-D�~���Ȩ`n;Y��/��G��&6�J@+�� ����}��Rw�./�O����ϸ��Yn�2Ɍ���G?�>p@p���O+f�<��<X�#�q/���Cmd��Z�O�g�-�ٮ�������GNn�~���QC���=��>�7��*�W�3&U>���bx�c������� J�,U�G�8�=��;��o��<'N�n���/�z >̛�;����L���'�m^���>m�+��/�tF�Vt���M��bRl�@����y�c9J&T�TKw�V���x�ɸ:���,D�DBc]d1�Yi�<gߢF������1x�4�nQ�NUB�Tu�b�-(a��d�_��h�>$� ��r[Pi��[��#;K�x��G07��sM����������&k�)�k���>��S��89%X�=���>�_�E<mU_��1��:3!k�KhQ�##�|+�<`�K1���l�ɣ����u�(�ȴ$�t3G9���B-�tTuOB����H�%f����z/R2nȬЭs���K���v�iUa0�OI�NP��nvfJk�h.oᴩMJ@��t)&�^�J�@JKߙ/�vJ�93�#Ö�/s��IH�.	�~�\9���Oq��l�U&s���P�+\�4�}u̬�;>|����ˠ�hI��g�/���J%�`���6�<s˲ »�%j�@��S/��y���rE�8��Z�����i�MO�(�g���C�5̑�7��$��zS##u��8s�:h�[���P²|�~��@�s���c��t��Gr��%��(�����E��ƅ�u ��%���s�k�5A�C ��6����kA��0Ė\-�l,�0�4�{ؾJ�N��V�/�h�;�<[)��z�e�rdZu�}�%h�	~V��r	�ܙ�$>�?���q��e��Y˒5:U���4��z}��]����f��z592nn^beh��٠E�ѷ��jR���I��=11�{�,RI^M/w�ʕ�3�
��(�l��P�jT���g=��K]�kmb�q�䮪ܢ#_>�*E�v�����xu�����]��:D���'���i��kޭ0��8r&��!;�׮E�87$_�]�g}���+=�k��ٕ�b�\�n��`m�����9���C�N��N����f]tk�E~Py~/ �G�p���h��
]�
E�%Ĉ(�{r5{����L���Yt*��M��g^+{��<��<��ig��[R}t+�ロr��J���둓|H�+E,1����{GD��
]�c�E��j~.��	6� ���l=ɕ�n^�[�e�eg�%:n)Ҁ��^��M���������|�q|�{���{f�i��Z��H%�PR��7����D�E/��s C����	�;h�$��j��f*�y��P{/�^ޅt8����°.��b}��W*�N�ߙT�{*�e�1�m2�_f��*kN��/\���Ǹy*����jx���Ѻ�%.�rYΗ,1��N�Q�t�<�S� A<`K��R3GDb��8�w�*� 2W�'D�f��	�}�����Vw�1P�"n|�[����Sthk�b"<O�c��L���?%�=Vd��%v��i\�u>ԦB�ɣ�@�)V�֘z��iL="I0����yd��,��������\��Ӣk�M`���-�о�I�Ԙ�0��V���ʋ��*�d���g�]�6B/��:h^��3��%��դ'���YfŰ�w�$邈��/�]Yj �͏��ZZ���2WH�c�?�f�����h(w0�:����a����Orw�@*>	[�K��Rt'��HX�Ac�?3�fs`Z�.>��cq�&�9f�	*V�4vp�^�Ҵ����Y�7����>h�� �쥷^��09Hwye��{�bőF���\�C��|�uCm���5�$"/#&���Ȱ��$cDR݂K��� [��x'/t���ut���Bil����\�P�;6�oEYx��|Jo��
����@�9D�[�8�" �Rz��į/���k�f=�?3zP�=o	�>����z���J�j��V�A\�k�t:�Cޒ@���bD��`����Y���\�,{�y��!��}S�O2d<b9q:j{Y��*=��A˱�Z��}f�#7D &+��xw�^_�/I{{0	�5�5�X�ʳ&���+E�Հx��\�iUm(���F�S��R'=S���'jH�s_���_H���<������܂��[{�w�d�{��ʂe��bʙ�#M��ж�wB;��]����-�/R#׭�V�&�2�ԳS��n��w�f�h�R�)���,:�	)��f�L�(�f_sF��S]�uvf�Ńj�Y�yQ�	p��!|�<��m�֓? �����a��E� ��[��>\��Ks0$�u���O�*��FE҆�/ޣ��<���y�7H[{%Lg�0f��e��!�j�a�H�Wj����?��J�?4��%G���W�"�"��Rmu�O�g/�P�q���̬֎�����Ri���[ܰ�S@�+��jA�׺i����6�xS���e9��ia�3����j���[H��L$!'����a�9=R�U`����"�;EJ�mI�������#j[gO�IJ'�79����0P�G���v��v�I����m���Wm���	��������:-:<�(�H�����I�m��c��|��� K)�H7��ʉ�У �V&�W"Q2ٞf��ɘ����_ބ�ҩ#��'��A
w��	{ 3���1��G+e�k��~Te��j��xp"=��us��i�{B�O�FH�k�e�j?���%�$٢������o���(;�T<f֤��BhT��(��_�ˮ��O]���k���l�j�_�tA!��2�����J[gA8H8������_�V$�I��c���?�`S=�������Rn�j��N�?�[��ՙx�� ��C!l����!�>	f�p2�dc��� ֍=]���PL���ë!v�X����ј�܏R#����S�L)��cݓ����"���tN� 2�x�IR�8�Եٻ�:�s�D7�+_����Q�!_p��9��d�̸��К%�����>��a�Fj#(~-3%�vGw_�A��Zb�n�U���X��r���}0؈H�ͣR"�8��$(<������N�<������� 0�55�� �4h={���tp�"e�	��냤�(���v�cr� ɌNr�E@4R^Yg��Gt��sK��O���8څOhOK��\0CkGa�	nվQ�ϻ�;PQ��f[T���B�h#�C�o�z��2�S'{4�#��4��ϰ���XlxVHYEB    bf14     c60�y�N�	��	���?���<%,F,�Y�!+�����o�?�8e���b%��#��2U��
!BdX�D�>��L@��*��nAPC��a�*�-�c�+&^R=������㨠$��J#����N+���*�=x&�qxG���7	Ef�j���k��mr���Yz�D0G���{1n�wr��N 3Ӌu�����1�ԕ�*� ���4-NJ6�O�-P[Ty�+��(u�y�]�`9P�]|�����9�s�
��M�u�w������'j��.]`:o�E�u�u�@��$�H�����%�\rdڲ���DM�ߪT	x��w��$�t)���x�.��5l"�����~	���Օ�{ǒ[��3��ɲ��Vu�/��)>����#�����RC�"�K�	|��+�i�fj�|F��}�a�0�k��?�a��T2�S��
�tx,�[g��6�D>U�l-�^��4uv�jk̼�E����m#�vcO�� ���h�>I�$���H���јu�f ���̍���/J��Q(0��s���1�n�Аk�S>�wk�mV��6�j9����M���YGTi����yq�@�诹�_/!�*hCz��u�=�#(/ΈE)�H�ӵ�/2�%���C��,�O���sR��%���:��C�5��g�*�6|�v���S�5�X�ڰ�.@pGF"� �P��VU���`��"�H4��_�:����S��-[�C��4n)�Rb	z�ܫqY�J=��8ڐI7鮲x��_�&��!������}��g�����ujS�z!����A��@�FX�M��Z�V�+���!�8��I�N�^����cd�)̝t���b�N*�'��[�G�<#F��������Yc~,�U�(p��5HdT�o@���pmG�t�fN+����Bw�M��!��2����O}�@�q�;j�j�����­�JfB���.ȳD��Y�*	&ZK'z����iE�1�շ,�����G�#f�r�R������Z=���܎�&=F(;��<H�N�Z]F-��gr|��7)��;:)~��R�,�s$�j8>���M�H��1���w�P��=�hv��瀋S�8�EF/�l�:@v�_S�-b���&Cݦ���5�u�tv�t�r�0d*�r([�������W��k�¼j����BGĨ��m�0�H��i��.�)ǅ=��}g��h�����Ȑ�
�#:���x�s�7N�o!��i���VtZ�#�KX�u*�c^\A!X }q�U����G>_��ƖvqU+�]kę8�m5��{9aŀ�)�[?��7����������FS�$�Kj<�u�!QSGѭL� v��<\ϖ�%f����sʔil�gf��0񀯝d�69�}�2B+��@�y�@�HB��	��h���?}�ͱ���� ��{�|?^�p��]��R�|2�o�>�c�t[����{pt�����>f����R]Lm���*3i*y��+9>  Gq�i������v�"ڮ�X�_���������x��+^?]�1���>�C;k�b�_����4T���%L�Ħ��j��}��=��P�v���@�� 9S���Ea�'+Z��|~�/Z�� N�,�)i�v�y���|ndR΋�@gY�C�eJ�za)�Z���i/��b~�PJ�ǔ-�C�;�Ԓ��B�u��(��3�U٬�sszh��:��%�kwF�����p������Ff�*y�#�hݳv�x�]��9�<��sgH �5M:�7k�~C�C�Fݏ�M�:E4���?�ߟ�.��q�>���s�;��c���l~h�(ط�G�tf��!Y�)pS � ��w��v���!�^e8�J�r�ʹ�?B��in��J�u@���6Ա;�aV^�w����^4��P�.��a9������sC'��IL5��5���l��kA(��{���� ����։�ͥ|�Ȃ�s�Lۤ��VN_,�`�"z�ʗw0�7^�ڕ��""	ZM�O�ί�/�����vS$h�|zf���9v13�xK׶r?#�k��w��t=;�� b�Bk�M����h��č]t���n2��O�J��CyD�-IMe\(���(������E�~��6�\�\����8Ҝ���TW�����1�4,��:P=���i��^�wӞ�O�D�\[�̎P�W#VD�u0�T��$5���?<�8�T�#><�5"����X���4n�4iVVM.v8��yd��>Lz�?�vp�~���(`�6*w�� ��os2D\�v��RK�J�2S��J���v��o�p[���kn(ߘ�tW�xس���699������xio�?U���6;if(��P��0���M�n�78�7���a[�DgË{��$�S�H�*ۯ����� ��= @~�Oʪƭ�Vj-�������G[b���+aݥ�>5E<��6)Hg�rWM6��nk�$6�k�ӗhs�&w�ܐ�n��>� w~5vӛ��C��lm#ςUh��n�Q;�U6���gD$:u��ܨ�����X���;�#G��%��` >��=�(��1�q��\F���;��|E �k:O��B��fA�P�f�ʢ���.p��v.�q�����b^i'9��8�Y?��	/+�rG^�?�����gIΦ�/AB��d��1��5�J�EQ�w�^ξI���2�����1ǧ��9瘝��~�?��ҽ��8Y�o��i������"!ճ���������V���|\�S�P�9Phl��[�$�4lzfd�'R16�T�?O�3Wd�\F�<�T����-8����H ��q\�Ꞝ'N�V<��"n�;|�씓Iꢉ�w��|79w�P« @��wM"�v�.ȶ�����Fڄ	m�3��#���R_Y{� ���l�^����z��Zܒڕ�8<�c���\o�۶�d���#s�$;}x�B7E�S�0�;XhZ;�
,�e�ed�^;?x�bp�3ͦ��o ��e��Ґ�w:�����Oeu[�fSP�/3���{N�Bq)���Z��yy�d`��̣Q�wn-�~|�q ��|5[BØ��k�{�qy�9"�bp�Fo ������3FN��$��J�-x��쾮�q$����!�m?J�������9 �H�