XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"��u���E~�x�!�P�n��2oT�c��uk��\.Vs�Ȯ*q&8&+���,v2Q�A�^�|�Н
�C�;l��[.>�I5O���o���5e?��.��ʹϿ\{�ؙ��{r`v���j2wH]&^#C]K�����I]*��� {fn�̕y���F,C�c����d*�?��:�D����Ň�S �U��������'[��Ȥ��;�τ	l��ܢ�$uݞ���$�)t�0�B/�e��݉��\ظa��b��[��/ �}gҚ��L��o3ܺ�/�W����Wr!�kXL"��d�^O
�%%�Y^����,]E��W��n�|gR)�xT��U�G���]�OC�Ҥ*,�S�n FHvE�s�AY���}�0 M�>}?T~�?�i$�uX�x��#��'��Z�W�Ԃ�����As�R�zm������<l,�]����`�enr�����8ɶ��ܗ����6�ǲ>��{�"/r#�� �r�VX,�.�( ���P�O��S�+�3P9�.S�^$(�,� 9COJ{
�iR�W_l&0����6-�=X,��D��2�u��F�ͩYV��餎��P�a�� {<�2a���^S���/A�#`k��!��HU]˱��]�&F٩�͋�4_2C
H��E&�<�f	�0s���;�!��Ќ�_A^��H���"(Q���U���!���C��i��~s?�w)p��Q��U��D����=j�^�*��'�XlxVHYEB    29da     af0�D��|V�fY�]�v��+ f��d���S���F�30��R�T��R���B���%�-�8Gj��V�߀ۆ8�	�&
�S����q��z����nA.��J�]��m\�k�y"3u��=lz�r%VJ�q���V�w=^�)j�(�@�,�i� ���?����������E�7�8"����VJ� 4�c��Z��G� �.)%M#�e�Y��K��%"�C	��|͏��~�e��\�2��/l�<��s��g�n�����͸Z3��|5%��(AĴJ��|Ya��|����Akn"οm�M+�W���.�g��s�ХM�ߌӄ��^-������Ѳ����96^�S���=��#���E@ F<����;�Fq	Rhl>��g�A�feM��12�4>�w����i*o	�d���ĝ.�iR(X��_iY2(C�}�`mh�n��tF�$��.�h�">���zi��	�N�
q*2�M�ø�_�:#�v����)i��\nھZ4l�ư�=��ƂT�}s���tv3P�!��@�%�.QmOV:�yX�[&��=�XW�A�xt0$x�ƹ�'!���5��3�^�����dMElT]�*�h�ǵ�~��Vy��?w劲X�^<�#�W�y�<���O㌇�}ґgP-���Z;�oSb�$I���|1: ���zDlC��)���a�X(#镳FRߣ)ɔE,w;�n�z��e���$I)�|��}�R�:��/�-�}�0�b��잱z@��:�,�h�2�����NJ]o:��X��w�M�\e|��Z�ݮ��K�is^�� �O��~�k��~-��hG���& �����!aT�y��Y��	ƨ̑���P;ғ\���X����*�0p�Zg��$��!�F�%m&���!���q���$�����~u�k!�Z
���О��*��)%���F����>o�Q<���_�叫��٬�V��w�D;���&"���R�f�1C�n�zTG�0b��md.P]A'��׍�1%����T�"q��rg"�Ke��2�����G�n\��� ���`��R,j��-�0��)��^tJe_ɼ�������S�G*���y��L�˨[}�~��W����$�W�f��}�:������Ց��@i���+��K(��x�����\ w/�������~�����9�EcI��n���؈�A&��R�V �+"�7n���I�R�e$>,�S�`��݇�@��0A���dtA��&=�P$�������8�4ztm���A�PUG<e�,��0��Q��k���w���O���54t����#�N46��C��j�[��$Ƒ�T�`;08M*����Vv�v�0v�1�H���ɋFg΂�kS�Ty��1
�V2|9�Hp�ǰ�g���^p�¯w�S}��d�Pۈ&�4|��أF��5��\@�����۲�:���Gf��lm�6�I�7�F�n���~<��3%�ʞ�ɗ7h0�y�O����5����zZ�[�-��N��o[��c�Ҹ�B�B(47n3<�zu�rai �ǐL{�S��4G}V������Oru�x�}D$'5���������t�X�����@U�b��3�}�IlH5�����5Z�����7����i	>?�k�I�"��D�L�EE� �~Rtvg�E�S�Ŏ�p�s���NN�U2�Ju���!����YC���+�kT��jM0����@�;c��#�������Z���+�������ㆅ�O�3�g-��+b��fj�S�?\�
oFd_�m�-}6�Q�Ҕv1�oѥ�q0��J�5�=eAz�SwS H�e(uC��>�/�� 6:�>n��:$�ǟH��!�UO*i����r�8L;�	��+�jl��'J*6�JY��<G^���9��������M�)�B	�5�����I�ǔ��C� �=�GR�g����A��Q�Ͽ]��k�� �;�D��I�4;��ٽ3��$DS�Ռ�Q�~�����K����j��6}럦8"�9�¤�i��܌A�>$(�=�a�Q���8<V��N��3����ב��Dn��R��ja�J����6}d�R�Ž~��'�pFQ-��/��E��T����IT��W�0:8���%f�,$p�
��'�/�J�ѐ�:l���`�,���t���N��:<ui�QO\��a�|���%��Cx���ҭ��8u���ͯ���E��?��������D��/��plT*��p�ˑ8 `-)l��� �@�o��A�n2�������?�ԗ��z��-�����<��x�Fsi%�4O��8~�ξ�����t���WǾr�e�"�
��#��H�5�?�8���u쐻Y^q��z�Ӫ���)t;�<[����<&��NKCX �\'�z�s�/ߓ� J[&
Y��+{������hnj�� p���:Q�ჱ��ly	�8��O!�AdqƁZ�r]���iZ'8�X���Tꤾ�Pk^p�ƲT��{�L�=����_SS^�>ĸ�(֋�/���s>7-	^�Q�0�&>�[Rm|��'#�g{�"���]Ó��Å�y�*i3^��{����߶*��k��И���4���W�)�O 	�%��X��+�K,��O�À*Ц/_5�'bj�����W(3m�1�I�B{ S��Ӄ>/Z.)��]7 _a�J,I`r�6������C[J���R�lM)�O�U܊X�G$zǰ!����'rhFǠ&(