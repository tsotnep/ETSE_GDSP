XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��mx����&Æv���gYTT�0��,/�?��a)�b8Q�A�b%�E��!u�DU0�2�ܹ��
D�[����tb��v�yHa{[W����T9E'��l��;����}S*�rB�{�K� ��^h���|�cx~��4T���JP�˛�+�:�e%���9/�� A>�s��X��9\.7k@\F`K����rN;��.2n��iU�Ր�e8(�{�A?Ǎl�T�	�!�l���Q��V�_xB��}B<�=�=V�ϒ�vb�AM��Gq�I�F�:�,4��q��"����ٜ���%P}��8����ɹ��u��IdHz��C�����}�a���Q�>7��?ןa?���[��lx-��,�q۲'���F6n���)��]���hF�t_�y ���E�(y� �uw�&]�t��3�����i
�$���6���p�
T�P��?%Y�wwx�6jTwu��>��Q3U�H�SdK��TǱTSb�.���x)uV���j���L�����[�d�C�$��q���+�T]O�}�~n�V�Ys�qo&�����~1��8K���h.����Yl(Ij�2��s��X"�`�F.���b������������&�
i�؉�3i�/7�I6N�5f�������z{��L�e`���ڡ`�������:����8?4�������)ҕK��z7�?��6����f�7����h�L�٠�Y��sˡq�N����n4>�x�Y�uK,+�{��I�����XlxVHYEB    fa00    1f80C�U�������gh>\.��L7�$%�$'eD�NkT!oT��#�sV�`��[N�cF�����'��w�A�00� ��UC��Un�����[`� ��O��{֋:�� k�	;��K���^	��i��;�o�.f�Ը���UccI��I�qQ\1���.>j���1eQ~��{ ��e"����3�J�e��Q�
?@X���~<��w�T���� x0�N5;�3cyȋ9�� �-C����t4i��0^�3����?�q��;:�[��bw��o��)i�@�LJ~�t<�@Y!�/�a�g�S���"$����<v�����[z3��P׉8���jU:����g�M�s�~|�)��Ҫz�1���u&��j2��#mBe��S�=5_��Z����%wĮi^���v��4�X,ާ�W}����[�磊���:� 5>��k��md-�mo��(���vɸ��p�k>ཉ�h-�������TU<y)b�u���-�2D�%�����~���b�\��פw C��$*�L��sqsjm 	����2Ȼ�S���X�O3�za�������]�ɐ.J i�0�>x��>��X���*�R_?�ևEVT5R-��6m���m���uM�܋���Χ<�Jv�����mk&U\X�A6m��or������Ș
y�?����4��6i�r�5�q9�\֛��h
�F�&��㷂?L�׺1�d�E18={�!� Đ�N�Ì�	R3��I\��b��o�����G�$� ]�q��u���e�\��C�6��vh&m{d�N*���9�҈��V�|��x�����ބ_������_���<ܯM1v�3��Jk6�U�:)������p�l��Yz���Nvw<rc5�Ʌ��~�mnF��9��"Z��h'F`����nP�İpVrd�����M�:Av�r��gb����G���� ���~J���[Q7��,�X	KV5�0�"pX�@�;���7���@%@����~\hW���'�>�{o�<��h�R�_���h�n֮V?��e��B}� ����Q7*l��f���G�)�,?�v�I�?�6�>1m�rR�x*���MI���3-�ɪ�u��!����vE�eJ�ٻ��v��nc*�'yvkդ��q�Dr���<Ŋ槣/s��2>Y�� �¹�_ҡ �/�*��~�E�J ��9͇[�e�ٰT����{�N����ރB�d�r������VH `��c���%(�#	�3���X���x���`GY�t&t��Ɖ�,��B�!s�oDC�r����2�]��lZ�N��Y,L؉W3ܤ��˟<����<B	r��x�uY6�ʞ�k�;�nX\�@ݎ��|)'})�K$��s��'FVE3i���U��&��I�`�3�j	_>���Y����ة������,Q�v�rV]�k�nY����Mj��]�Q�+�Ai1�^�M8k�~��b�{�k�w��En�W��V~��\<BO
�H"u�MRCIa2/��|$N����(���G��%37��*-�n���k|�@H�����Qd��+D7����*��٪��x����L)>�+�$�#� ���WQ6�j�P݈	���w
]��sөS���aOBh�<pԕ/������)�a�E�M��+�B�x�֨����ֿ"E�G.Y��9.bd@��q|7,2;ҜD`"z�jMn'�uH���x_��k2�:���_p���������G���V����f�N9#2Ac�%�ϴ�S���Mʂ�\x�V$�9�y��\���p)�n���~9�u=w��s��8&�����&�ZX�D���'�U�~!w�:�t��9�5��W��|Y1m�K��af��jR$_���%O����ᄳ@��*�� ���U]�2��U�/'/Ԛ�0~�n���1���9��f��b�N7 8nR�{3[`��3�y�F�z��wƣZ�\�+�7J('��>�X]�0Hqf,s���H�Cv��R����9�8�_�ա�hr}A(��ݐf��%q���Oz�!�Is��⑲`=0���	1�p�4���$X_j���^��$�KT8<�Ϟu(�����H'�|1@�b��f9Rt�f
4'��)���!j�i.B8m�& ��PoǢ��,:���͈d1���n�5d�-����o�g�ն�����K�ԗY�>	^D���1P �:,�v�v�fk���hq�V��ո�R���*��˙s`ɳ��F��:���޾l� ��q��@��*v�����XuURy)Wi,���Ӧ��X���+8�E���K�Ŷ�>��Q�0)�PP.3����b���WG�R�Y5a5��js�S��=!�n'���&�ËUD+ _�C�a0&鴁��r���
��|���������B�n�����g&H�F���f����T��$<��F�H�yPw�۬Ě��A���g�q�cҀ�����He���2�Ј@�e!�|Q��!���/�ڟV������qԢ���������Xy�\��t8��y;z�d..Nz��f	{�D�<��EN�h��Ļ���y�Y?���q G��+z���D�w<r��:�n|�,̀�z G	�m��O^Ӑ��YQ'(�{��S�M�"l����U�l\��ϟ',1��G@9jcC6K^����s���3O ��J�>u�-^J6A�ź���m��1�B)I��i'�����^~K��=��!6��s�|�sƯ�!��� c�ο٣�A�]��Wd��^2�=A�aO�Zؓ8[s���wL��5���z�*p�ks�Ӗ����YLf�X0/m�\Zπ�P�=Pێ��xɕf��.��)�cû�JD�Z�ZǍm4Cᴢ�tfRu#Ţ�Up�φI�~B�)�܂����wڛ<�8E�r�p1¤���a��:�^ �<�?j�;��o��&���Ͽ�j)4l���@&|�h�M;İ>� ��0/]r������r�u�[��a�CVB]O��꼗Ќ�6G������������L =���_�P�oƆ��
E�����b����b~Dd����
�Z�>�ȵ��Ȏj>ԧ�Bv%v�W��5u���2w��iȚF;QZy�+�Id��
9��U�_�
6�ˉ����d�pf����a�ŷG�h6���W������!�	��/BU����̔k�۶~�t��oM�>���?��T�={��[T�)\E���������#�Cֈ��X�qT�b�H'Z:���Y�]@[0Xj��	�:��{B`h�"���)m�����bK�^F��L����9Cw=�~rG쓜��^Z���f�pN�iG6Ty�껵v1�����w{\;��2]�^�������*4��W��Ay��g5,}��4nRO�v`�l!r����zq��aD=5�F����	�Id�FP��Ց���G������/?��%^��%V�y��ܐ��@%H�����U�{��ː�Ь��e-4(���l2��wgR�.�UCٝJ`��02��$iA^lμ����Xnդ}��������4�5����d��D8���+ !�{5c�&/nj�����%BɿXO)���ہi��M ��:�ے��;<r�#�m����X�؅&P�L�Ta5|�Aᑢ����(�u������������r��6W�hP�x����QYB*�d�k+�<K�p���g�Yx?�i�l�(��|�� ?V�}w9������RN��<�:�!;�Y+u�X��&	'(~��H��yjt��B��?���|�z�H��{=Z�)�Ν����m��1<o�"�AM�����jOu�;�q	ٹ5������b.=�|MT����-�{��h��a]� �cV�9�>�M������c��=���Y%�l�q�]����))↔���x���4 2����|b^b�2J�Y��}�t�V��wV/��×Ayj뜙�ж4/�nD���位G��f���uF��\���d���ϖv>�������>
���}#kp�X؜����W@Ѡ�9��]�,�[,>��u�0b�� ��j��ύ�js���+���H.�rI�
W����(A�(A����7����{ yA(B��jl�<W���qQ9�B�)���Jbj��Հ����\�\��O�$ll2�bҵ���,��o�Em��gj?
��*�2�s�CK뺦�W�)I�j�C�q?gФ_����[����V�����%�	҅L@Iy� ��d��fƿD�?����Q�s��W	��u��S'��j�\�����sd�{\�%
0Zw�M�.[H�����*N���אP��M[�Q���J��}^�2��z�����x����<�&}���`\$���t���*�2/mx� V��xS5�HOZ�nU'q
�<W\�&raf����r��e��(J�������z���.�����b�t���_��3�N#�� K�٬,񹫓c쯧I�F�i;'������S�����g'}�SH(%I�����x��/���f�-�b��LQE��N`�0�&��S8���b뱋���Pvͼ�dja"����ZN�ٳ���!��_��t�9��5L�ƀ�(F,j8��%��Hh�f�d�$&�0� u��&���4�� � B����ێ�3~�<ʤ���=�g�lc��W�g&ddk�!�E al�]Q{ν�!�縕��H��I��PĔm�f%�MG�FPEc�A��y6J:�Z�$���i�z��5b:�	ꏛ�[p�8��ƍ�5���&@Pw�iW�L8\��(S��&�5���Ey �.o��G�q���ُ[)A�6��V|� w�)���B,����9v�Z;�O7�/�'��iq
��s��u(�rJ���k&Ň���ء���H�8��U��};4/�7 iI_����� ӌh1I�6���|��FO�!��T���!w-��`�p�2���_�F&ɗ`�yю?�[�����>�v�Iv�z��NՊ�o����C�˼�����+D$5����)��C���b%�]/�  ��T�K���0�A9�4�-��+aY3K�8��\]e�����~%���V��k�m�ʏ�A�.7=�Zߕ:no���7)��G(W �3h����)��v����n��qJpJZ�޼E�Bd���&&��!��+3����l>r5<K0���y�@�̗�xMD@��^�Y��i�>Y��jC�]�`��`��	�3T�U�r&��l�XU}[�@ۡ�m�(Sy5��HC�|p�� �=U��fbس�[�qn�ܯy�	CUb/�(���p�D�y��zOT�)������\ds�ڻ����G�Y�]�"���GW�kAcP��g�  �g�����'�ٷ��:	#X�Ml3�$a�3����&UU)a#�OW¼�k����t����Ө����qCۄ�N��}�Ք�mۮp��-z�x,�IX@�.Cx�x�� Py�l�5Y�X���p�}t-S�ނ]^���ʫ����Pc��ɞzG��P��)�&d��f�������r�Ѡ���_` �B��V��ɚa�qQ��Xf�lv��Q�*i�3Lʴ+�e�~������cA;�����4[����no���#�[��` �:gʩ��	�h����ڊ�#���ئq�;<N�?�\����1N���D֓�U�{�~��y*�׹����o�Aj�hD�D�vwsQ#�D�.S6gC���ao>0�qy���'!�͊�X²����A;-��ۺg�G�00���wH`Y��ԥ�t"&hփ�{���C��×�l\+M�ӋHa�w҄���ڌ�λ�D4�t����obu�ؐ��\�J�4��n0T����0FeppJ��ʛ�	g81K�)*�9�əs7�	���g�56#��RqR���+����Q��fc5�NΉ[���G��4�R�Ja�r��@=_dg��*��@ӌ����Hʮj�>K��'u�K��r<uP�!���#!����o�	��V���C�]&)�Hz�':�]>G� �^9��Z�N�'���l�F���bd���X������1K��+�-�
��{�֓���QAFa�y��ǼV��z���)���
'��E�h��V��Ff���X���P
.��C{�:��� r|��:j�z쇉��{J�j ���s��,y$�#��>��p@�涿����[��ڊ~s���ޕN�fs�z%�w�hpx́g�ȉ���+�$��6w��e�I �f���J�K��"S���Զ+~�O��?��?9���1���P��
G���ll��+���?1�f�T����ak��8����\�D2��[��#5�\V䝠�"�tVB/����~��R��Ys��h��$�ă:����YW��\9���!����N�1S/����8�<����^��%�-bB,C�����.�x!��x=��شA���/�}`����>�׵�2vʤYg��Tu$�I}��j�ZS�r�M����Fy	�d\(J|:���+#��u�M/�eC�:g5�Ե�B�����#W�Z�'�үh#����~��B���`��<t���;wہ�Y�4�Y����Io���wJ�c����=�����v������6xU�Z]!��_.h0g'����c���;t�����`�4���6�(\Q�`v���zkvE���k��Ze��@���
��4�����s��7)�u�T|���N�E�^��RYO��#8:��۸&S�[?W�f�/�)��e��7 E�������X�|�l}�\����ɨ��@�#N�'wC1<�F�!&q�M��*$G/=rVK-���t���j8�LO!�G~�������9��r,�fj��le�y+�n��|�S?�L�RP3����-@�C�؀�[�K�:���SP�<z���@1&��g��m�>Q	��Y��Ƥ]mg�m)�L&����5J�}0ɥZ5�"�� �7���RdH1Q��mR#�T��5T��ovɱG�m$�$�h�J6�y��'/�օ4M|w�o�$m'��a6j��4����v��5��+5_e଑��_��Ϫ�Z�"�f�W5��p��[�ꁗܺ�)����&�gW\�=T�Q�t�TQt½�3Q(��o��V1��q�b�qJS�a����'Dy%��"�*��?��+���P��o�x>���LI~���e<�=�ںvk6���d]%\}��7�w㠌�V��%��^���WRpƼrָ���%'DEN�q�g8ߠ��v�2m��qyZ�gs���;��e�0$C"C?��9�����q-&yϋ	C%��Yr��M���.��g+[&Cm�]�!s�`	���F�"��ڱa�; P�"H[PK&3���c�h��sOڠ�n��[i�4�y��=��v����Y窂ӶaM��XH�s���rT�*�Wވ��p���c{6U�ʹ�_�����ù��(̟j������UY��v�\�S��BƤۡs���oFP�d�F��D ���R����U]U��~��%A�b�D����%�O�����!ʼ���}J'�~�D{��EP�i�|]K��L)���P�b3�G���4=z�+)�;j�\�y�@Bt�t`U�/��@ �����SP^_��T�Ղ��<��Rgqd__K��}7�$%G�~�ʄ�evƩJO<�P
�7dͲ�X/v���{����PP�;��F}�rR�?d�v�nA��3�s��U36��"/�9���L��CR`{����ۤw�`v{'�=�Tg��޺5UgO�C��(��Pۅx�Y).t�Z��]��}���vѥn �63ilG
�+ծ��ַ�$�_��ا�8� n�K�Z��$c�>r�����a�A�I�3ig*�:V����M]�,���o����Ɯ� lj801����(���R��Z�t�?�����v���z�XlxVHYEB    fa00    10c0+��L8���������>TtbeB+����5X���8������e��$��bTo�]�"�5�F�
 /��3�m~��1P u�	�h�)L}�s��Q;�6����B{m��eS�i�� �iG7}37���&�俐w��pz�Z^_����a��������6��Jq�&u���8�P2����� �T57Rm'��.�]򟃟z�#N���z�1�̔`_����`��^Pbx0�Zw��5�^ޡ-*ޣj�d'�e���N��"o(c����$�����x&$�\o���O�d=&�(�M�Ә��^��F�8Q��C�|?K���K�^�y��u�\|���^ݔ����N\�!��( ����j9Jf+e�, 쯑�թ��'Ƨ�X0���� �S�'zwpw��㨔����Í-����AE�6�}ű(�s��+1S�=�S{e�v��4����R�b����u��I��Q�ֳ��	.��V%��T�x���9����Ҟ㟏��
Bs4���z�?�k�,�(;�f�5�|�ʹ��z����y�CW�- Ͼ����GGtg�c^OIB�ʮߴʚ������Ƙ�qh�݁YxVL�W�d�Uh��×�8(q]����gB
U�WG�~R(`x�xd�W���Vk��QU�V��jb�ac�~��;���Y�MCb��lXJH���_B��������B]p�3XR�YZB�M�^I����|��zЀ�R��k���{'���r��@R��
Di���8�Y��?���VP�����ꡙl5�_���(���$�#�!�BVJ~p����vT��r��]o#4�cO���߰�4ܒ�׬���g�i�l�	�R	��u�PI4yғ�c����ȹ�Jw�8찱7>��η�C&,�zg����<0F�������M��w�%����)���L�a�'hex����m��(�x���E��]�r{roSv�NA+/��#σ,��1#s��I�S&�������iz;k�i�i_�M� 6��ƾ�J#�ڢF�����r����i B,�/������H�u�in�2d`n'����g����iQ\g�&�2��G��g_�w��ß�p�m
�\ IL�'㘩�oҝ�Ƿbe�xU�p�D@g��\��R3�˸
'+6��NW��n�J�����I��J$�f���[�����qW�Fqq�f���Y�LF�+3,8��t���+uEy��Q��E+T5�0E�U8����0c�	ٙ��	v_��2��o��ja���D �j�ǔ�wЪM�{����V?��X�����}�ˉY�*��fUKjY|�N�@y��^S$���9)�У.WP���ī63L��y}D�4f������g]��>d��C�R���B*b0��˦>�4�4"��hs�b*M^�I�����V��	�F����M>\+�x�1@����#��s�P����e�3��Tw�N.�����UQ�&t�.B(��:���7_���w�hw�|�*M�B��(Q��z����M{���舢x
6YEm�i�*�I�hh�}r~�������O�ߚ�2�r93U�of�Q+��NY��z~Lh�kyR=�di�(Xv7^�����3pJnexMۘ�RSo?O���
�.���j�V� W�i��~�@UN���\HC��HRCt�x'���39���6+. ����S�,�5Z6]�����s�"�l]z�����
?�~�P�ݜ��)S�A��/�����F�f�v^u �)�P�n1����3�<Ĉ�G$�O{���3q�,}I�6���G�/��t}+u
A��e[�q�KC_W �.��0xv��Yے<��E#�n��h���F� ���%���[��,Ii�-��*�@qz�m�V�#�ζ'��
��P4�d{����~8�����D֛��:w��G��3���;���J#�Qҡ	�`'��-&�/Հ�+d��6�t�Y�G�x������Q��[�:�JP�+��Mk6��[P�ɴ��)��ɴQ��v���&�W��¤kD$��?(#L��ߠ(��^�⿘W� 4-�Π�����:�jք����(�m74#/��5O�${.�Z+��L���ϧ+�꫙P��]��MP��7t�p3	s���TU�Ġ!�1:1�sa�k<�=��cb�|l��{�"�^�������:X�1;ݦ��0�˳?�-64(U�Wy�N84A;"]k<��bf���L��9}�����[�HP_4��63�(Z�Uz&rd� �C$A����h�"���>?$�̃%X�O�|⡠Ktha,J���pə��u1��a'�B̝8����d|�D3��zG�q��%E��Qwɫy��P�
�z�d[{Q/{a�1!R�`�#g5yj:-���EJUxg�-~+�Xi��k�gGm�f0Ȩ/I27��>�}�Z�����9�7�Z~���L2ѡ�s���w5��ݴ�iO�c������;�*p�]K��?9ت��ܙ%Uo~�����ݰ�nq��_������,Vc}~�j�ҩL�g5�wWп7͗�	3�О6����\�e]�ly[z;'eO	+�D�Wi�P�'�.�dZ���9:���OEf=�		�,}|q
�OO�v;�+��,0�hQ�Q��1G�.*�ӄb�t�OL��{W`B��V*t���A��ud�
��Ec�J�B����Jƺ�#m'+;�$���P�v��(.0K�<Td��G�4+zZ�X\�y��f[�X���O].�z�!<�=֕sx�9)�ٛ��*�g�][ '*K:P&�a���맗{o�
����i�Ꞽ��ۉ��hɇ�'׋�"��ZDz�������V�6����%�����/*�T�&���GN�9�h�K|���#Q!B*,���̴ZڕDCS���M@fq�7��̇Q��J���!#�g���H���|���[|z*�;�do��F��<&##L������O,��b�,#I�$�y������6�;��S���)�����b>i[�vFGVC���:�d�7�?պ����A�a����Q����Tz���6�K��&|v�<.<e�hC��,�&��1^��r݃�#�b+l;�͔�>ON����񫵠��>j��;��d���.1�S^�l+b �&0Ɲ�	����hɇ�3�k\!��EB����d���O.���'���sÝ���/�	"ZO��d}w/C!�$�YII�����x��H	��q0aV㾤�ݶr��2�Ş���r�!a�^����P���?my�O 7��\�b�ت�f��"��?�w��%%����'����+��]SOȚ���tm���Y�q�eњi2F��f��; eT�E�N�h��k���	��"�ޝjHr�/���� �y�rx* ��c�Xic�]'s��E���h"��)f�������c��2W�t�D<����7Q� �s���
TV�`�+��"�06�hj��e�=~l���8z�7���S���j�Q1�Ա�9�[�a^��Go���x����6ѐ���&#7!�,�ą�JB�8����6��?2���,]k�T.���/~�jh����V|��s_�X�/�iHR��G�ݔ�; ����/�S�Ib2΀|c�CT(�c3�qb��N���;�Q���r=/i Vڮ%(<���4u
c�ix��=�⮶�Z��yo�=��Qn�5X��>{6���_:fM�#hW[X;����2�����ƫi�y:��d�Zdp�~�ݐ���s�ep�g���d\��v��Di��N1,��ygA���{� �tc��U�@��hOZ�N!�G��ets�Y����5�������3G�	O=�l����"�+02DX�.��(㸻٪���8�}ǀt[R����k�?�+a�%�*(3�y
4���>����#���B�K�t�łt�����j�q�)��#�$����
�=57�Q y��6�Z�P`�{�Q> -ni/�R{�\���@^��ꨧ�B3 x�6B4��L�i����2�f�%��턬���9�U}>�?PP �ø��ӜJ[��Z�U��b�Zs�z�h"�$N����m#%f;�DZV��&����}	`�?5�rn�$�տn�f5l�|uz���}��G�ݤ�m�g������V��ZA5�B����O
I��у]��=<��Y�aX|���|�:sC���,H�;�R
��ɽ���2��g-��XlxVHYEB    fa00    1140W�[��lY]tXk�4h'K2-�0*�!�P
���h�@��Ɇ�$�9��*_^����[a��Ӽ��iE ����}�?��&(����p��+�O�k$L�2$�$
���u�?uan� !�KX�Ȩ�}���X�R�D4څ�5�a6g^�����5�2�e��I�#^hn�gh<���B�2�����<oQ�"��٪<�XӁ�R��~�FU���q��
Җ��F�s����_������+E�%Ӷ��cr�����n���o�5�ɹU�=X�!�."<zU���-����4��n��ҝ~=�|g����(��E9Y ����b�Ք&�ξCiŗM������P0)���ӽ��J�r�.�bVð���c��\U�MMwZΐ�ES�}ǲ��e2�����ʒ�ծ���{e=Db*��!���q[`/�;��m�kGB���:k(�҆9�q��r ��?:�PA��G�ё����-tG�ӷ?����	 LD���F��Ћ�`��k\��{z-fL�%xw�E�lU�U�c��J����b�[�q����l��9.@��1�ee/]dC�a�*����&���$��U���	3�1�v�@�PT	S'�ɱʼ�b����b[����2*��6��N=�~��1Z�Rb��I��^՟EO�Žȝj��F��7�괟�5�������U��[̒���c�v;�P^Z|�S�m���H6_�Zn/JC�˽���j�7**V$�L��2N��?�A��Fc�<�݃�
��q+��a��^k�&<F�Fb�H1Ғ��4�P�R�4�l'd>�z�K;ͤ��� ��+�?�,���e'R�3�y�`�����u^5�[2������2�fEY]4~��7�����gOF$���J@h�j���ui����;�U0$��>���(!|�������	��R">��!C9���I��4 �v[�10+ŨO�j 2��G8�3�ƍ��e��ԩٴ���19`��-�����Bp@�������ٴkHB"��I��.Ĺ��6e���p}��sgIϛ��[���~��� �f��{Ft�Dw[i.��.0(���
��z��p0q�7�;������!ϧ�:���ꛋ��t|A���5)Wl��۽�[NKi�����;,WSX�gk�  Qfl��CM�%�(*ž�tX���Ћ������C�����+.�%W
���ĞQ;~��a74<ԕ�#T�+�Ǌ�a0t�����ޓ �x5C�.JTK��0�!�h3]+~"��V�Lci�����
[���Mָ�M���}�C�/��H�⑹E�5m�C�R�j�tm����5���v>�镐�����9�h�j}��P���©�@�3T֍�-���� U�d:J4;���l���*�NȄ��q���Q'+��W0��uLQ+��e�0��m��U;�AyN�Դ�e9��Y>����'/p��S�
0�j8&�/��
��b��u�L��k�Ӧ28�
���wc�)sW�i��/�����=�q��q�3ßY��u� �B��c������Ļ�~jMcW�(���
A����}�N�m�q�Im-%}+?�䞁Vw�R(�n0�
�ke�61H� ?��B��:�RuZp|�j$�\	i�+lҁ�N!ي�L�*��b�������AW��3�V�9��[Q.�hr9Q#�ab��[<�#}�b�^��D���AL�V+�=�B���Td0nQ�k�)�P\?B���cRP�/N�O�VE����������2�1��R4Mv��\v����d�X��jJ3U|	;��L�_�s��~�a�Lr8TÃ�!�%V2-:��)�Ŧ�k�ןD�@�i���G 4��U�dP�����~�d�nYG���D���mb�ji��N������T������z������@�Z'pf�1��_&����)a(�����4�l˛��C��/2u������{|bZ��"����\��,J��U<b�W1ql�ߟ�9[侸�]IPA��0r��@S0<^�m�ż��(��}x0J�����8�m�[�w��W��X��_b])s#�g��b�M��w9���.�m�\)6� ..��_�N'-��p%9�M<�T�7!y��JLY����B�:�1¤��B�����!��΀�q&�w��a��}P:	͎WWʊ�\���v����t�y�m��v�<˳�r����{{����s�,bX�U���| M�$���ʡ���*���}U�E��{� KNe����*�E�$���c������V�9}�_h=P
*��S�����j��)�q�w;�o�����+��4�;��%��8Z9��C�I�x�M?��l�{���>A ��k��9����}��м][�+�8��Kԉ|��H;Z����껲�%faM�r���/a��9� E���bv4�V���D��$9(�F��DI|�v����B���^�oy�ztNK�.�1��V�Q/�i�Og�:���?�M�R��^�q�mU�o�p���Q�D�'�E�Fѐ���7��V���Ȇ��U�+e���^kI|���z��候�H�5+�"��/9}IZ��O�Y�p�˔j]��?�R'X?�o��a~3�� (�<�� f\�ˍ�2Vv���p����&Ƴ$����O�%��e�M8��U����Ҩ[�i�ד^��J�t1��ٰ:��dD����"��Yq�R��4�\&s����/<�?����ح.Щ�/���;qWNv.��i���Ŧ�S�-%�~^�K@(#N��hmO-����?�ޟ��X5����
L~F�"�_;hR���P\���F�S��Л.mx�f�PC�L�1�{0�Yǽ+&��1�0���{L�I�����#�����d�d׊�`��+��`e���,�r�STQ4O�x9��B洧��;��W{�Cr��u��sd��$�?��x4D��J"^s�QZrB6�g�7��AW�ZR{��n4Y[S�jq5��}	����P�!�ȳ�)hՒ��l��q�bF<��E����ԫl�Aъ�Vw��&� �����9���WFQզ���a����ۚ��C�@ G��Ib5�禳�J�P�u�S'�E ��{P�ҫk_�k~���ԣ�n�ȥY:������8�ɽ.��36����!�k�p��#��4�h�h]D�
a,�ʏ@K�����5����	L�BYe�^�d�Ҟ^�c��:��7�Mz�v��\(z����}�J���w���s����;6�,j�a���j��p"�:�w3���b���C�-ru�[Z�dY"1���1�yk:�&�� �Љ٬�d���>+��aݕ-�I�p�a����>��a򆡵u�����?dV������0ii@�~�6���m���Z�L�)uRʮ��2s��=�ϮĀ����<�f/GΫ��W	�QEBtt��Y�����D8���Q�:�ㄻ�\\&�m�/߅�����[S�����j�{{�Z����2,� �����y�W���ic�_�9��	�DF8Kɪye��b6 �!�~~{���+x0�^��}�zcj��·�s�X����**M�緩+���|��ZBcx}6ZA9�� $J�B�ꐨ�J��_�$��qkdp��Wj�>���u+/0�p#���oh?�<=����D�C��EP=����!���w.k2+k�y��������M��]%m�X�Щ�y���)���C��u��s4[�(N��Bt9]�p�7r枣���%������]��X#sm��Q��ѽbL��E:���pr�>=�G�*f/�>o���ɡl�=36�L<P'@�Ο�7ey��d�*x��:�7���P˼�n;ve�wSH��+Q���^�B&p���0�q��هջO��΀�υ�W���Iф'�p�Q�H�y6ݹ�M�T4�ui�hQ��B�n]�ʶ8S��F��h+`�,.R@#�p��Ðװ@��p�����yd�o���ͫr���9g1d֕n��$<���7:Wn ����1Ru�>?[�I�g 4/3)�5UH9u��jE|�\^ā��޵�� � ��y���4�er�td^��9�L�\?�9SR��E_���9���@u������:�za����Q���W�#|tuv�Q�o����3E%��B
��\mYyدӫ�n$�]E��V��\1�|���\��-��<x��g~�B�m%N����9�4�7A����?�
H��񡕹��ѻú/ `?8�
[F_��Ȯ�.��xi�&%�8e�xZ\�)�;xD�L�����}�`9�;QB�X9��d�[ B���}��h��O�	l�>$$XlxVHYEB    fa00    12e0�� �����p�8aH�����S��X��h��~��Q����m��;���[��vݳ{�H[��tmb�\�[�2W�r��ώ��a|-�2�:���K>�s�S��ex�2Cy�K�ܒ����r� �6#��C�m�*Oߒ*cX��P�r�I2�����vH��=��_�̗��(q�z 1yq؉l�,�8;�冹��N�J� �>/j�C8�/��Ǻ*��zm���<5��
%�9��e�X��.��D���&�B�K�o���f��]X>�՟V����I6���H�`Cꁡ�gx58Ej$�M I�(���Ð������4�W36&��ﲽ+�o�c][DH��]ӣ�}N�S���r6��@�9j����Jt)&�b�ڰ�{���D_M��G�Z���ϗY�c$����j��R��@��X�@�s�?��Y�(�+���w�(�*n:K��5��GL�Z+�};&ɀqm5L}���^��s�@Rʃ(=fC��/ý�rɂ��x�s�r��fŞp�	{��T<az|R#��k[��w��j0�
���Z�WY}���mLrf̈�@3��	�?@A�ʍ�oB��ɦ�6X�sQ��ֿ���[���js[DpH0�89��l�t:�V�T��J(�&�z��t�����P&�:����x\A'�~�wCך�&v�����p�霑Ih{1 �] �%n�4|�/.�i�I[����fc�eo�}�S�,Ͻ�TH�`K���jFy#��0��a�\�����U��q���)'�2�R	UT�K� �E̘X��
ς��+��$'N��*���TR�����/��C�:D�{��:�[`������r��F+11J�5zV��,��F-�������H�+ ���!�Գ��Ax4� O�C[��B<ln��Ʉ{�\����V�=o�T\��Z/K�[�h��T�JvڹB�P)�#��̸,�����C׸��1u��$���?a@%됤�6ֺC2�?�vefeqDP���ϑ^����WF�2�K3�I,t5�ϖRG{0ML��{Ok󩡓�e[��$���OM��7��|
��� ��3�Е��3=d�s�8Vˆ�⿫�[j���Ļ�H��NnISCy�3��ڭE5-�?!�
�Ȕ��~���5����IP2u�<up���΀����pY�%>��;.m�6Ľ~��NJ���Zn���v�2
�f����0s��9�yk3��533���Q�x\Pǐԡ�DO$�*F�bl��}�z/cS��t����-Ҹ6'`ƥ���g�/P?Zl!��C؇��Ϯ�zY��3n�-̎+���6av���33���k��/��o�נ������W%�c�� d+��k�����׿v�R� |R����|���F�h(��S�����@�ɡ��o��RՐSb������ͧ��/ ?���鳒t���5g��D�@t̳��'�a���2�%�I��A|�T�K�k�WI�/ z�����U��2,�q�UE�诂*i���ړ��Է�� �6lU�ҕ9��������Lص��錢aa���쯶�͛zкRZ���0gPH�o��4,�N5��xe��2%��a��D�P�1S��j�[Հ��~�6�l�ؓ��f��V"�� �� *����/�,��%�!��Ȕ]k��_�=�3,?D �DD��[�X�����f�%^���1�[��lE�!D/ՄFDh./��L�q�׬�;�N6	+6�Ǌq��w�嚽e(<�e�����n�T�sg)(��L��͇��%������Tu�y͜F{���`u=��$&�B2��(����'^o�A����o����#oS���nWI�[Ng��B%w��ƨgF�lܽ�Q ���+$����q�6N@���������bir����A���G���K�+���5H�
]�]��i���h+�4+#�J����V(�.�\Q:0`��N4~�*K����X�$�,Jn��C���@����C�mN?��#0Q�5G8*0*�,?�^���|���:TfZ��6�i���Vq��W�0ps�O�bz��Bww�?�����>f�՞ :��3L�:��x�R�8a�����?VU��Yl�����''����3փ�0/�%��y'kYR WcmY�k���=���R�����3�f��6��f�A�e/)�0v&�ە���@�˯S��ל&g��S����U��4�"@�@��B2%�)�n�Th�\�Ŕ�b������#2{#������INhA��{GZ� Z>��sKl�7���Jq
���kc�%h��V��כ�� Q�1�W�����	�ZM��`n����nS��`�&�uX�Eͽa�K�B����&�����̕�S��h���Qu�g�����4R�C�
5u5;��I��3�tm� ���>>�>�U<�¼���N�W�tfB N��8s?��yت}���yUB��?����-u�$�q&^*�5}�\=Vv��]�ͩM��d�oX�b��dtu�� ����$|������)���׮��������D!�x�]ɜ�t��܉������圷٬U��l�z�_�'Zn��U��UG�Y����>����F��G"���ߝ��t��+�'��ɡ\y�"�?�k�E�8����}�v�L�p@�G`�_���`�&�@����;z���Vxu{���pD2'��h�0ˮ.G�[��=R!ę�l���y� N=�� �97p`zr7Eh�Œ�������n�e�����G7�H@A߷��[�D�"��v�: B?����坼Q�`6F���l�����"�;]���~��Pt��������n�v ����ϓ����Xw�֬�_K<�%�D����ѐ�T�OT���^� ��,_lg��TgFJxy�!���*��㊛�~��[C�[�ؘڙ�6S�.N��|Q��w+�MpCHy[��ya}���1��Z�"X�iㅊ���U�f�|\�A��G��/
A��d(�I<N�}�UQ�L����$p��G�#�2�  8�������(�����j=V5/����wb/��I�����r6$"�%��-�w���p2CΤ%A�3�\լ�;J� ���Ħ�:�vO�#���za�mD�u����x+Qhd�
��[}�)�[�Fb��mR�>�c���]��Jb	��W����'��l?6-$V+�p4_�q��Wn"8��Y���Uq�,������5<=��D�K],ZS�C�`{���	�B�8��F���<�o4��9}��ƚ�H8q#�����&�]���`���K��%����8C���@ B�=y�L9FXSx�[�|���!r힌�,�V]i�e�jt_�ſ�[&�2�k�iG�Y��с@�C��6e
ַ��=4�,����k��y%u�
s|�h�P�R��Α� ��{+Z	�7E�_e\p��MP����#_���nX���K/����P��)�)�h�rŜ�]����W*'h�]�I;+n�J���B�C �SP�u����0���g7���U�lv�\� �P]�E] T���s����x���Hp�Z�u������Y�i�mt�����g)1"���SG��b^9g���Z��M�"ڪmkz�(@�$>�k��M=H�KXv%o��\�5M
ϲ�%Mw�efV����ݟDvM�����Ф=�C ;A�Ysh�Z`��A<�n�u��Ë�Pe70jjU�>]�~�!s 7�;<�P��:�	MX��O�����������9By���~�E-�K4�1ɷ�4�6/��`�y���w?��;���QrĀ��|�(w��R X!ѵ�9��x?���!O� �� �+T��)�R;�𔴇[�s�Q�P�S		�v���pyZr%ӣ1��II�����X���lv���稿�z���U-{�q��1ۉYlqR�Wg�(�W��>'.wH��q@-X���5�	�7~���֩#�,j�dl*�sD���~UG���<���J2����)C-�]�b���P6fy;G���~��Wq�t�L�wrr`7��B����f�ϧ���,��o�'����^���	�eF���pA�9&�j���.��+&%k��5�H�<U��&{z��ʤɟ��Ya+Ż�/��*��338V[�b�z3�|�S<��0m��G�P�����!N0�|_����=�[apP��fq%� L��I����5�#�4d�-G��h��Zl���rE��ID�G*¼}U c�4���ĠNt��`�����X,ĕ��i�W\����A��lyQڃ]��.�4���Q�Y�y�a�Dg�d&�yf%��5��[��ۏ~]�=*8#��f��ϊ×�����)v9/�u 	�q)�
<c֯M21D8�)oyj�bD����E*n9J�[�}�>�a{̓{��
�����}�]�
T�).~�J�O�� ����1�Z��ʪ<|Wb��(w�b�������3�c�̂��t;��g^~�Zv3�dx�1b��ISmBw�iO�q�*Y�a�n��G�����[��DAM��4_���8�S�9.D8$�oө����ʱgR��B~�
|dWdM�9M�0�����9���L�����@���{"(B�DD��jqg���M�C�U�b:��v�����?CM�sѵ'.�zy?��{�����mN�M�,�X�@E��E��'��6�XlxVHYEB    fa00     f50�|4�`�� �x~���3F�aMA��VQqD���H�;>�1샲�<PƐ����@c�rK����[�L[{��.!��	��'�*Ar��X�*J= �#9sk���r ���>�ɘ�H$��T&8�C?wN����D��W((gK4�PoQ�����B�ũ겜�������x�m��2\����}&C���RV��s�E�BP��)���I�fںXD#�h����+�Ɵ/K�
8�X`����s��4�@a�n�y��T \�2�	�6�dYQ�,�M�1ԧ��Z5:%�vJ?�Ӯ�B�&�*�?�I�.�`d��A
�Np!gt�}ܙ��Zn[�熇���V��\tt�nv$*ɥ�;	k4�d�ی����da_3��eu��k�Vk�����A[�5B0�i_ia�!C�|�b�YC*!���J[�=�:�<H��>�����1�$roz�gV[�u����U�ݴ{0E�o䆚XH�YF	��l#Ƚ�~-׭N��z"`��H��J��(n���@�`\�R�.�M�*l^L_l�A�F��ӤE����r�Swؕ���A��x�S���p�d���ms��㊜0�w�c�!	7�l�&���#�oZ�^*�5�WK>�{J8T���E7I�{�r�'RZ�4p��b"H+�e�@F;'&�jQ�K0T��A?M���Z�����.���8�\<r�A	�#o_�	�3G#K�8�Z}S���=��j�F�خ4�v!���S8re�8܃r�r���|��4��>�͊�nKa�:}'�%�M����p�a�!�wMzrך�,��{g��b���:)*jf2	<��H��6���Qu�Cٽ���ڸL����\���p��A-t�̹��5��H�vN?��))ة�S����+7�t%�[�r��� Ώ���g}�L�?e����!�)�Bd�KK�΍'8T>@U]��T����@H�n�r�l���Y�g�E�<��\?�=�C���>X�#�#��R!1�t.�>����`�s/)��7��(	�.7-����46u�	(��ґL��>�[�H��8�Uƻ%ѷ
Ȥ�����'���X�B�r�]6���`�j�vf�v�f�H���Y]bO����>� ��C�)��o�7�mG��LT�ĢIҰ&	��2��d3~�Iź��b�� oa}�'3���ꃙ�4\npsz�/��&�V��7v+f#��T��t�:�UTYl�>gŝ�C���ܟ�r���3O��U�������n�t_j)\(�̓�����sB��zO0�.>\�=h�mm_���������s�gH�;��f�X���Rջ=����WySI���輓���P�럤1�� ���}|�r��]}�V��qf�Q��TI/�#�5<�|�H��,���IA�1��G����^�қN��8����ʈ�BX�F5�u 9�Kz�� ^��2ݧE�)2�"����60t^J##ڼ�j��<���C�o��r#X jƔ��p�G��.���eyNN9E��̓����O+�@�mW����[����AУS�b�0��3�g�,l7����/G�庎�a]�l#�-��l7����z��~#K���+WrC�^�����}��c�6��E�3�&>����4Z�qD* "��tp2-�sn-\Y��ΊHS���.B�e`���e��{&�+n��5ȰW���]b��c	���K+�͈�H�H᫏[P�ldiS>�+���s��D�fw1��ձx�=;k��Q?�4]fF���}���=��d����y�,bڢ������0����*!bw\�4 �*�O��t�)��j��U�>w�5t�������>������7�l�?c�={�h׺'��[.ݞ��Yض�rՒ����)�!�p���T���3FJV���R�:��#�>LzP��q�!��۵l�, �JG�������bM9%�����J���,QU���F�A�V���h�X��8=��}d�^����ʍ���Ab`�M���;i�>zLlH7���5���?�ZG�z�,���ym��eD��G�8�ݚ�����M�{ŊbuK�}�b$(�6 tz-WR�H�C�q�Z�3[�A��S2߳���ᾋ�J�!��,eM���*䷡&���7�8p^��}9�{v��WLM�L�W�j��hq@��T��q)�~}����弘�c4���������s�?0���1Y�����]:��FJ�x�3fNXUN�F�j&�|:���p��u6����l0��폱��B�$$馚^�yRu�/�o��,�h���?[�Fg�_���5SD%�k�����LI�Ix� Iy@�h`a�J�}�,�9広����Ep"�g�l�(���IU��y�Gs�t����C��-��2QJ糩��Cl�f�����4V����2�X�!N�DK�F}3���
{坏��#M�E��{�A�?�&C�2U���I�0;�d�.@������M2ڇtH�1^~�"��~�
0���:[A �0��G�ʧf�{(N}t~�.;���E�ѕ�1��p�����?�f�ŏB:Hj&{�8��d`s^���X��'����L+�;�2�%JYfrQ�\�t�O������&�7!sg�5��v�j��=��dT����s�W�Z�[N���miW�d|�#O	n<�iT:��+���7���Y�c����r����<\3y������;�����}n��y#va0Ӫ�oJ1�eΜ��?NqUD��iqXy�:Rd�p����|`��	��έZ�j���!F*m�wk�JV]��"�Tc��_�CWA�>�LJz�a�?`�B������Q(-��$�u3v�"�}�d�����L��		���J�N[�(G�������K�ċT��W�_KĽ������ ���u��F��c%A��v��Ts�U�p
{�?� ��m��K��Z�j���2\�����������rI��z����_�E�Џp"��YkSB��=���U#~]�q;e���2�`OPp������k@���{�����u��9<1��[( ����'4�)��c=+���.�5[Q��n�39�-f�v,� �ab*�^���/gTȝi;g��R�����/���*i�O�Lt�z��8ڒ�������I29���M���{��0�ry8��h%��!OH�X�Z_��Ӊf���t�Ejb֢B�d��<���9��]�tJ�_�$T�"]1�S�I=D<�Fc�lo�u\�����<+�	5��-n����d"�t6���5+_��J &wU5}�����p#���i�kbNpvX�`T��C�ʧ`H|N�R����5�q�:��*pG��KI:Dtk�j�	�x��fV]���w��I`7!�e+��1��Y����w`F�x�c�5�}@�[O��F�mg�QMg2�+��B�l*�5��,햫K���Ǘ��b�V7O��c)�`o-;��«���p�����\-4�eR��*�y:��j�|�/����`�]j
�4l�
��?@�W���q2��NHQ��˻�;$+�*|C���^O�a� [Ǒ�*��,Y����m��F!�(rq2Vœ#�?��%�?Ӂ
|�hP�P���K�f�{�dI��-Q����,�{�1p�;��!���D<�iG�*��ɐ���a�M)P��P��^�Y���sy�x�V�9w��:��<�4����
V�B��٫%��+��b!cU
�����T���˳ߢ��VV��l7��S��y�Н7���-���m�JU�Oѣ�W|�)e��ji��$�_�������`�m�'�N=<��?X"Zr���W�N;��k���.����aNx�@E+�h��j|����t�
�Q^,�8��W����%��k���Y���ne�mXlxVHYEB    7273     5606���`�=��
p�b#��>���x_J��!����^$��� ��]�;l�
�7d͙g�ӂ��%�:ԟ�N2�����u�QV��#�B�1��iVۑz�Tp�7���2~; ���K�t��R����.=(����x�b�I�,,���/�����ou�#v]���G��S���ט)��]��kY�{(>����H�g�"*��!k�Ư�%@Hg�5yA���}��.��
ۚdm�i|��cҔ޺�3�}άl�P���𣨎����ʔ�Ţ�˞���Ҫ�?�y� vO�T�g0(�Lov�.��4Mx��B�9�"4�EG�[@��Q���7%��z���u)�*�������j������4ai.aa��^WN(P��'_q�z�W�tڦj�������-����kRr��Xi�2�4Vn(P��>)��|����s9�du�Ly��?<ϊW��������&�5!�0�I�d��Bu�|��!`oKE���<�i"�?e�&͟���CV���x��^����8���vi?���1�^�ɼ�_�pD#g��ְ�"ia��㔺=w�h��w��Lש�U���`f,�62$p�E�zGP�(�耫�WT[[mNe+���wK�ϐ;�)Z�~���H�R�UbWM._)N'��F#,,�|���f|�d�c?V8^^�#0U�!$�O=�n���M�IO��9J�C*��q����"㝜"R�����7���ݙ���%8>�j�H6���Cv����v���R�1�</�a�`�@�4�F+�f:.T�9�/��W�5�^Su����ll�;d$�GpQQ
��ۀ5�����E�O�^ο������pD���D%�`w~�+��o��,��y�v�8QF�v���L�p�^뼟oJ;A�t�P�x[�r����cgi�k�uRK�}��lq��YK��$���b�G�"�TZ�38�U�y`B<�/�A��'s�TU���ق&
�$��Y �cY�V���}�F5� ��4����Զ*����J!GW�%��5�_�ɡU	��==�Gw���P���Ob��~�G�#/�q�q�z�S<�J�C��y	���L|�ϛ��~P�O;��U��P��##iR��)v�iu7Cc�����G7��훐���N�vs�B-(a��$#S!t]���ׅe������w*�M�0�:���0R����ЪlsI��ł���Нu�S#�r����s��-�4����㦔/^Ŭ^�+�����XM'?��>|체�/;$܎Q�>��-�Ǆ����[����e���2�fI��Z��*&�L
E�3a��\���~ʪ�����(�b)��#"�Xj��Y�c�;/�,�uAte����4��e�A0���x���_V�5�x��_