XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�o
��M��*A�DY�x���%�p-Cwҋ0`l^щ �Þm�Rm(5B��X����?��*�n
��IO�/K�F˔�l���V��Qa��FC���7\i������C��q�eK%y�۳���H��.M�A=%���%�R=���ւ�Xҧ�t?.%Rq�DX�!�;�����X�s>�5T�M.��Ӳ?o�����Xx��~Y�V����9�@�Ms�Iχ�<u��+���+���e���3p-T��:�aq�Eo��Sw�;����m���H2iw�4�fm� ��Q]�d%!Ϳ?�i��εu��6��-�[�3��A�٢���#�1�f��g�q�nZ�k�ݎ�A�lUx�@O+[x��,���ߚ���-��0��ڎ�)3{�p��{5�Ӎ�"����Q��q4�X{	,�3+!�|��'k�N�92�,��%Q �%������Ĩ��$��Ԫ���e�<T��������i�� ��?:-�G�'��$�����y�v�ec0�`�/�m{jG�*���N�I����:����xPȥ��$]��k=؄��.�*/�xv)g���n���_^�a<�A̤�L<��O��D�jd��Ѹ���5 ����Q�@@*A��u&H�_^.���aK�b_�s�j��7�,�3�ϋԆ9P��C�G$2WXgk����Œe+�Z)Vp�lT�[�-�����'�j�<՝pb LW�ĝ����->�)�Q��g:��uJձԐ��

��iǏt$;
[	�QW�2XlxVHYEB    fa00    1950�eo�x����c��f'�|D��XV�׫�0^�D�d��Q��DH� kK��}��`>/X��%}H0����n��l����!'��Q�e�1��_lD���AJ'��ن��*j�:IH�^�^�e�b@'�!`����>�A�*���ҔC�s�I�ѪĪ"!u%��?�Z�t���҇�]�ze�.O�Uq!_8S�7���g�e�2��p������&U'�yYE�E�h2��C)3�w묋��^`5�ĸWި�
>��~vK��E8$�*��R����T���j�(�>�-sC˜D�ZV�G���4�������z�\Q4���Lb��7.��C���H�IA+�7�(�f�	}�q���@��0o3���������b���-���������/�\��B�r_gK�1�}��;Zה6;{���E�(QJ􋵢,h�`������M�p4����9_OuR����G.�?�f��,�4`��\qN�4�8#�:�7`����}���権-�d�w�`كX:�d�@z��1HTL�_��EG��>�ɡ��}=����g���x�x�6�t)�Ν�?���d��x�(8��!8&Ծ�F0���7��aj �xBbY$��F@��7fy�a %��Y�j�{gb���th��)2ج�N���AR���;	i�V�~6t�=R���][��Q��w�	�M�����>���aiO�a[�q�~� ���ҟ���9b�uD�
���Bv&0�|��UZS14��V�Xt'4�߸�j��} Y�xk�4]<��!�Ʉc�S��`��0�}O9.��q�o��}�2�p�	鍜}4qo���-gs�f��L�>�xM0�ީS7�j��W5�,��֍�"��2�)Q3sND��\pȬ�	�'1d�'��-\1HL���x���Λ$C�}u���9�c3gJ�e�Ag��A���鷚ļ�vJ"��U��ۑzW��������1��Oo�۬Ҳv$PN(W'7aY�O�(��a�9]��@�5�}����Q��S����������u]L��~O ?A�8W&G��F��n��%�S�=�O�ԥ�b^����������Y1;i2z����#����Ӆ��6���շ�Rz�h�]����=�ƪ�f8�9��W�7ɲ�B��9Tq�C���#�G���p�q��)poS
/�>�į~/���|-J�q]7�n@�v� ���������V�GXĵ�n���6�u�;�L����jɺ�r���*�=���<����*G�A;��[��>�n��[����`�,�%d.� ����BY�!��j����h4$����-Zû�r����nAV?E�ה� ��y�Y"Il�ʯ�n�Syy�2���NL���[���8Bn��O����m�o���z���J��Z��ڹܠ�a;u�k��Y�:�b�SS5O+��'��</�zm!Y��&�Q����c�m���j}��YXE���0��ݓU��' .l)(N�H��XAD(�^�񗀲 @I]���H��^h�8���#z�-� �j�d��@j����?��S��j�����#BD5��?�u��ǟ���۸�N� ���s��h`%�{#R:����v�h����C1~,]��ஏ�,�r�U�����gEz�`���n��?���G.n%Dm?�X�/�a�*BtH��ҽӊ�m$> 0e,��GFI��Ó,�ޡ����Y��E=��U(u����nP��s�<���MU��s�<�N<s�`��[L�����!7g R�U@9�P%�xQ���H���7�*vGkNn�}] �Fh��'c��j�����HW"�l�&���Y�Eż0���Hg�%�9�^����l=r�JW����mM���M�$�����.$_L�1�
A���6����3Q{km�&i{��դn3�:m�q�������Ua]�'Fn�+)w�Y�i��"ls/!ԧ��ܒ|y{�Z��^YгMV��|�p*��,SO��Ӗ�|���@��e���R���XV�Ga�5<�}�{s�ށ4S���I
�<����d��{lcj�.�mW4�P��Ŝr>pp�"p��,���g)����0ؕÉr:V[۝�,����N0"ڷcN�,�2U(������Q�wL�w`���@�Fs����Z�'e����{����=�skx�dQ)�R7V�r	`���#���|X>=�d��u�Tn�.�8��/�T�_iOv;����e����!#�Xu\�Ö�{^�w�]�׳YH�.��IϾ	cp�Ͻ1y���OB��쿈�<�Z��o�#x	���G����S�,�0;m��E�!�����	?@~מo;�0 ׾�L��c��mQ�F���]�����7���B��Ň�"����. l /�F�dw34��3��.���L��2z�E��6��FYk���l�o���;���6�����������D����o���3F�Hޑ��Wm��JЎ��Fܗ��\��P�4b�E���\������^�\�L��(8�-�u�ހ��@ZO'�叝�V�U���-�6��r�
G� D��pAθ��IVgT����*𸪂�p���Tg�t�����Ɇ�A!Yo5?��b&�f*�F)�Lgm��a�Q��
��[�:�:�O:���c~7��P��D�jJpO��f�a��R��'0C��c%9��4����1ox3)��J��	5��\��^��wĐe�����`�"w�R^׹�CNLJ��{ n�g�<9:j�u`�v5z;����t�5E\\Ev���)~�d�th�?��8f7�E8����;в6���W0i�� �3����-K�~�B��d�_;
H󦢸�;�V�*��>U�A�^E)�����vC/��`�j��<E��utH.�Φ�'����(&Z���B�]�I��}oc�Z�GH�
p!E���RCC�lſaH�.��ȏ��~Պc~��t�;�����1����3p@�ꯣ��ۿ����-�
���z�C"����%s}�	Xʣh�J[�������Ŗ��u���%_X2����� ��Tx��R(����_>]h+�M,��;��4��W�Y�1&m]A8���l������ת�� M��fL̻c�%cf��T8����;��(	�������𛝚��l�Št���n������%���/7�Ɩ�Z'���i^W�	�_�vT1>�e��@n�D�V	�ʶRD� �2������g:��s"=�u��x��Qe�}J���*{)�g
POk��ȸb;���E��_s@7���߁��2�-�I�ʜ���f�d8
=��h�#OF��fh�5ů�W����s�V���}>�$$�� ����φ�OZ������,͂�v�`��d)�evH�Qt��H�L�3�]}�A}�I^Z�j؍e���w�Z�э $�6��pEF��ܡ|e���;�%�w}�����R_:�'�[t�L�(`.hJ��9�y��i�y���Za��pS|�� �[yb������f�Xr�{�,�,���Q��?=
�f��D�]P�-Zۑ�saƨ���G��mC�Õ�#�oM0�m�l�W�l��t<A~e���DT�v�d�� �~):#5�:���G����.�s�|c�?� ����v���S4���R�g>�
���R:fIQ�v��u^Y�j�F��Uf�޺qF33�jٔy�C7�;�g�u%��xb���V!C�����6~O����C]�3Asq��	�9-��O��j.�5!n��:���X�4��A0K�~�7<�L�R���p��)
�����
�&���l�����N/�-�	��䛕P���m2�`r�=�i^!�N�y�뚙[�`����o��K���D�{�D�"Y6����P���_(Ю��w�s
��.88��Q�ۖV�B���>@�����N�t�K�rJ��dK��˓�^��V�,��`l�F�8�r�hc����kBw|#�꽏�m�ƛ`4"�"��7��_�u�.l���ݗ�:���*ÝFX[0=u+��K�Ʒ%]�i�ʆS��+T<V���R��%DN �)���W����3h��;԰U�"��aɡ�u�8����e�8+�$L,89��>Q����+�%��s�Q��R
f~�r��u�|��^X�� �Ì#���������D�M�0��(eaW����x)G��6T�j:u�|(
����������d����p�ǜ�V#_�X��	��?kv�>̋U�;�k�X^�u��+@vdu�C����(�f��Y�7�6�c���%�p�T�Q4eɞ�[7��~[�}�����Ճ̒e�%����I�a��<�[چA<�l1+R�B�De�r�$��u�+*\�Q��2���C#O~<����� �W��Ш��{!o��!�C2�܎����.M���C��9R�x�jMz��#�b����B���QRA[SeP�9������4��U_S8|���#U��S��@@�u��.�=���b�
u�2�,~3l�50>w�{�M2�h�s���-/��Yy�|�FN��yp�ҝ�x��Ԫ.�CK-)����[	���Z��+I��.⿽��QT0���T��i!UD���=ŏ�j{�T�F��X#���mp����4�]��5�(�+��`�Fu���Wxc�?�iT�#6�`:��Z ڥ�7@�]�$;}B����H�O�Ίl�O~p�L]�$�k��sϥ�pbt4l���Ə�붎�~�8e1\DHn<��P�J9����:��]8�J��wX��h�D3-^�zI��{T�)���^V !{��?U���az�jn� (�̬��Kd<��+�LV*�	��ʻ3���GL�)����������Pqs���u�39C��.����Ȩ\E9+�7��2���]&FaZ
�j2>�͚?�����,�@�U-W��-h
����i��d�
Zi���A�Mvp4�)�MP�G��@�UTa��r ��P$h��֤[�ꡱ�56)�(m�n5q]A*6q����T�S�K`��)*yY	^�F~�r��=0�Zg��i�F� YZ�{��6�5)�-2����p�+h/���i��Ɖ�Y����#)���)
t��Q��\n~!Ǩ0f�f�@ݏ8�fk��.L��@Ԁ���	Z�],n9����/
(@=��GH�J��<2�f5H��9ҏs���~�,�:*��cr�汜`tA:�f=�L�8���9k�Am>"��V��=���3;1J�K	��=�ZB5�ãV�iP�|H�S��K>�F�����~«��Aj�@��0�9ɂ�D����s��5�rf�̗{8�RQ:�E��
���������� ���h�w���ө|�ao��l��U��#��@�ﬆ�8	��u��H�b��SE�g��^%�!�Q��w�)�"r��8�}��LZ�EՖڨ;�>>���[����{�v=w�D�KQ�g�.?���5�M��M�Sx�L �g�	xn�@��/��Q�v$��tP`W�#�ű;ݟH=*y����|��C/6�uap�ɏ�פ�!�s)=̬��Omg��/"@�A��� ����:2���0�Mn��\���[���5Q	�܊t9^~l�I)n�f%~!���w�sK~Ӯà(��8g��'	���Q���$�k�v����˕o�I�6*?b�}l�`J�BN�b�u�9s�
"#�3�^C+�|�M���K(����aE�UQ
c��Q&���N&t�$+��5b���.���X��s؛��$7߀31��*f��"����G�v�����s�t�}=�$�R�q�b�V��U꾏_^��fnK���,ol͹��������I���/�{x&��l�-��pܪ�4��$��^����$�9| ��
k����0�?K���G������+�봍�6Q.6N�M��/����χ�g�`�\�V]9H�~�7�F�,��d�k~fj�[4KB=�fb����
���2���^�>� s��4��*9p��'������r|���������2�w&G�|L�0�� JS��b�bW�}�&��&
�����!���t�t�cO�P.�[�����w��)�)]<�� �i�� ��R6N��M��*��)2ٚ�T�
8��VN�����Dz��v�2yiKD�� ��Fi}c��R��zd,:���Ô���'b�?�q�]ޡ�ǳ��q��́��?,�i46�<&	�{>��ĭ�`��*�,45m�`~񙄒� �t�y�c�LG���t_	�r>�[�Rfc5�>����Gke�l\��{o�����O@��H���!k}U �O��ݨ�=��n9��I╞�'�9�]$~��v���j*����|;*�0i����'˥�r�H""��ۀ��ӎ��/FB��@?c*�@�gɇa��l��귏��(��-��I���.�N���~"^��2XlxVHYEB    fa00     700|L��*�~��y�<e?�y���v�D�z�*WN�(n��!�/�H�	�/�M�f9���� ��~��W&R����T:̧mRFe"�΂��ߦB�ܡy��"re���6���"C��	�pCֳۯ4.I65�+V��k.�~�8��Mµ���{����Ҡ�.Ψಭ>�m�
���^U������WH� y�k]l@G ����r���DW��,��KRt��q�M˄o�1��/�=@%���ZC�('�����ZH!�峱5m㻈��b��b��&��e^�Iڋ�ʔ�]����b\��H�A�c�-���~8笻u���L���B"����_�#,5&�J�db�P��mJ|=+g%C.����
Έ�����$߁҈��<|R��|uS�f��:�#̡��4��5�ʣTO�@u(���.�q�Yҟ+�o��E0;�Ov3���7;2n��:�hxC�2<v����[�u�EvQ��Qu4LRE��9���.Kqp�r'3tϚzP��!�]�O�I)*b�tVF��o��N�O~Ng�Ӳ2=L�]��q��@����lv�Y�l�&� S��*�-�S5����ȵ*�Œ-#M��Ӧ�5=��.�{����T�c�����Վ��C���ut9�D�q)�m߶V4����c��h"���2��"�>@�i^�eO,"�l,��9�� Y��<�q&h�t��.��^�;�)��N���V���u�)M���5��i��0�����g�eօ����9S!��z��	c��<{ ŶMH����@B-�D=�7ԫR�k��U��lm�S���J���?�;�d�ed�I�aCB�=q��>Ϝa�{��9�o:���Z/�3i0m6O�Q��3u�d��ߴ �7��L�P����ㅲ(q�R�a��ԣ=��֓oy2 !l�m��^V���	 �5Z�&��$�>����@U�J�O��`�3��a՞I lr�D��;S�:ׁ�9�Y��P��G�Θ�նƜ����F\�J�i����f�@��t�|���ҼT��%�C����k��5�xy�W�-4EI��bOW4|
���C���;�]�V�nS�&����Ϡ�ŚO�3����IGqN���CՆ�W0E��qhlŜ��G����py��O>�Y0v���ʾ��T��TF��m|�7(m<����98(^p1����:u�2[*gSG��B��"!L�{��)�P{^����A������&����<w�������{.������Y�)���������+g��haRPg\�7�j$�o����3_K�g��	�t��Ͻ�*�2ǙvP��Cmfj�/Bᐝ�ȇ��Pww"��W=F,���y��w#�[a\\Q��aS.c��J��`�M�.�=�s�am��a&�N'�h�����"�@���i�+9S+`'�t��S�z-5�j��T�(4s��[W%�#���3�j�\�����U%�K�Wi+�?J����{��]>Q�yc��rt"��������ۂ�vdӭ��A�x�1��t�s��h�S~f��w&8ͣ���(��j�-%n�dB�觰`Ӹ�4���6>(_��@xr�b��(#�4��L��&��<�d�R���;����V훹j�Pۭ�C���R�&xmg�u'ī�@���<Moq���z2�KБE�lV�Cm"�E�o�w\0a��46�y"�z������}�^��\qGPz�j"
����;��?3����2<2�An4�z�DXlxVHYEB    77da     a60"�F��o�n:d�-PЅ��Sx�_�D��PsY�%Y�ڂ�0&%�������B�� ?����]�����dP�&9q�.Z�.Plĩ">8@�>HKY�;ծ�m�������Y����o�0,�8�)9Y; g�c�$J�$���젢�ɂ"�<��h�W�cg�<$q���f7|##��0-�3�'�-����"P4䖳��_*���Tm��J����j�ș��A���^®?b��ǡ7�zB�i�����*���f��?�����U�"�#	�iq�D�1]�>�g�s��z�xBG��+Z� !�l���*�^�_�m�ap��2ª�<U2?�!sR�޴px����� �nNt�Ф6fVX�!-ծ-���H������Q��f�1��>|T��x��zۑ8�Q�
�J���A�<��=ϰ �4��x��]i�`R̀��U��cyv�'Bޠ��L��C;���ht��w!Y׻vՐ9x9?��O��Jg!p��)�8h۹	)�O�uR����Q�1FOuX3�P��c��D>b��Ջ=h���w�𠕂�k�=�ut�����2��`��d��y�]�;	��x��!���vK��짊��M0�<q�����)@�,����χ�Rm�W]��!�P�%�0ğU���U�?�?�ė�������A����}�W^�F�갰w1������3��V5`�s�������;�Ե�LF�E,(�71�'>����hrߦ�X19"�4	�s��GG���f9m����?�'�<-g���i�y)�R�t��c���J��;r�"�� Sc���Ou�U��N�I���N�k���%�|B�[��LL�r��U|5�(8[Y�r��$��H\�V�*��dB�$����R#ߑ����x������{߶�`��z�]ؔcv+�N�w�X<$X��½�ˢڑ�$�+��K�!*Q1��a�]��m0�Q�����h�x���5��J�È���]9YG�`�ڡ@��e�颷yf�v�(& ��n�ml��E���X�Z
��3� Hć_��s�N[��c��ww����!n���*`��l�4�nի��uQh��?�NT�����A�'3���t��uA6Cq��{�I�a�jݽo�lw���2��ɍbnX�(���"jm$������=�	�>0�Zt�7���bL(�J V���$�LL�LK7"oϓF��F�����z�!	��䃉R`h�����xE(�24A�%@�AQX̓B>�\��g��:�f�N���ay���
�S�J'Qtm�/��^���L2cȑ�^�{V�u|�m��.!Md��ޕcą(A���P�V_�ػ#�v���O�5�&���0d^�{���^*o�Ot��75E3�k�*�!�h�]�z�z��a K�m![an���iy�.e��w�?au@L����h�*�q��^~� N��B`I�����!���-o�ٕ[��{Nx`���F���o���.dC:!��=�b^χ��ʶ	���Nn��%��J�5T;|u-֬?S^U"lX9
7�Q	���LJ��X�@�_b ����P0�M��!��71�i�j(���ӯiJBl��A�wD
�d��u.5�*	;�I��31r��WBb
�	���i`�a�@�%w�p���?նPU�g�P[G<.��&�#��C�� �$�OE�5���!x#e)�l <�ܝ��\���r�H�֓���Y�k�s�Չm��v+��\��7��BcQ��������L��7u�4��_խ��ށU2p]��-�5u�-a��BR<�4`<Q3w��ξ��O �h&Rǜ[����o�������Ŷ�E�!u;9"~m���	ġT�i٭�����	(��4�u��%O��d�Z�}\�	�y��V���^i.$�2v��U2݃:�=��%�x6�O�_ؑu�P-��ۃxCZ��c�)��)����!om3����a���:����m.K!�YaG}W�`��4|��})���PA:S��Cj.������aU:3��с�/T�3��B������WɫVK�*3�Q?{ٗD��SR��=H](�t�&�aؕ�����2� v9c�h�>p���{F>��Cp����XX��H��P~� ��˝�1tu�s����]K�O%�!1$��9ۻ��)���|ߴ�\W���� 3�N�MF���=τ��gp����F�1��'��+�I����g(w�	b˅U��Lc������X���TJ�������q<��|]��#��\B�lJH�?5���ǹ��]�G��z���H�{��vn����	ŗ�)`8x�jw�fxN�]������+���ۃ{Ώ��6l��C��g!X���1U�u�ݞ��L�A�|�.ɰ�Gh���ϲ
lxf������W]ȳ�}� �v��[D��N�畏��A;9��o:�B�_^���CgQ)��u���0V����5���5�t3U���p&�� ��p�]B�����q�$��#Ժ-+*������ �GD����������`�����L�״��.���p�oe����3S_���\ ���B{�k7�>\�V�S��*$Л��1��;��b<;^��i$��\���V><��I@7c��#�:Hpn��