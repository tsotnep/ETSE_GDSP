XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t��bm�o�)[TV7�v�!�����j{�.�D��?�Ŭ ����8�A�^1�H\����rg�I�ߕ���N\=�m,U��Z-Ŏi��:�|�>�"���x�PrU5���˸&��}�����W�L��s �GE^	��G]s����lsv��:o�6��E����I�����0�tﰑ>����ql�뙅f4�>a�a�ץXR瘰d��j���Z���~M�u�e,�Ju�D�d�@�����	9Ș�S�۫C�~�]�a݊��D������_��JS���+�	R��J����s�;�0�^�,��t/�EYf�y���LA�.���h�d#�멸���!N������p8�x�FJ �@��D���O��+jH�V��?'�� ��o?���t�K� ��^"ѯ�~�_��M��Ɖ]D�u]s�h3W�}����sxyB�2BS�'��IG��8D�ٶ�V�M��CV���������,wBO�	%�vo©���eT�.{U���2���v��'թ�My�M�B�_�HA�%������iD����I,q���N�@�,����kȦ�#ܑ$w�{ֈDh�݌n��EFe~�$48>�匂q���h(�K��ER�R�������0U�NuW(B_qy���D��OQ�^�?�f_���G9�
E\�8������Z�1���;�m��0خ���u2�n奒I�u�H;�W��n���?ן�y��[N=�R=�@�(J]u��:6�3�XlxVHYEB    b8a6    1ac0س
F�v�ݬ#  ֡�ž(12�����is������]a8�7'[?��3�W�hD�;�"�T]��m��P)^8![�U�@����9��y3\I��¿����M��;廫M�����jm	c�PuR�ZFq��ٹ�$��"܂���Zs%쬡R��D"$���G�֩�u����am�@Eړ&�Ť�?��3�K9,];M���7�-i{7gL���?H]/\���{K�� �pN�x�lݞm��瘎H�c��K,Ikh���=��֠�q��o�(F'�60;�$��H8c��d@�D�ޑPP����l���7��oQ���
J]���A}0�k�9D�:�����	W�EB0�P�|��z�ʹ2޻T�5i��O�}�沦  ?�p�z�0{n�𶵭hd��-<��&k!;��x����7�G^�v"�x)����h+�[�e�&s�݄]���j�\��O�ot@�7��T��Sϕ����b��(�prb�Y��~mBE/N����e��e���A��A��+U�M��6VC��b�#��A:D��V��o���d�m�bԖ!C���)�KBUP(������ٱ	�[�Ӕ%���)�L(��z2��c;|r8����w<�I�]^00�T,��ΤPb�:GVB���y�-�FA��0�L̏�<"�>�v]L��Z���:��8A��K?�A=�n<TR�&��(���M|?�k�\�ӟb���'�ر��&��@渤G�"�)R��
�&����f;�ԭ���L�|�����.uD�l�����Q-�����x�zI��q5#�Z��w��U�y��6H-� ��@�b0p<�����)��LrYs����9+�;A�$�u#��r���ÎD�	?�PV�c��D՟Z�$���O�|�U�Z�"�;_��p�bS �s����6�2qO:������ع�D#�H�06�0x�-~�T�>�(�<���>	��0��a�����ϲ��=��Ԗ�Ưց��^�?�y�� �=�$4-DXRg�C�{:�9G��&R�lg2����?���%@����Gy!�y_&=�x��:6:��~�r����~�-��`0χlR̹�D�Pw�refX+�dа�{B�;� �m���Ԇ���,���H���M���1x��}��}����nԷ���Ě'q	��� �T:�|�.ަ�=|@2ޯD���V�#C%N�CE���4�2pyy�>JjMe=�?QU���-�����B��;��mO���'5�8o���4]��
��ȡ�~}����7�a�)�geu���s
.�n���W;+��ZS�jf��x����R��ŪR�� ��-��.|r- ���F����^��h='����K�.g�ε���=�5ou�v;����L�(���'��&�}��諻��T��%�I�z<�������br&�_����~��O,QN�׀�7�%�w�!��g�6C�q饚��@�?tG_����v_��Δ�ep�UO����!<��C��+�,q8,����ޒ�O	���u�G^���&g�x�/�5��v>���4���?�7Ws����,Q!.F4�SF��T�$��:)wP.u@6� ഏ��k��հIpWG��H5,�>=&J
�[#;�.�+��zo��@Gu�����lPsD ��-�� ��3�8`�~�<����s�ڍT�_�!Z��F$n�;#�O�j�|L�,�	���&ހ�ӱ�R(˅�Q����,]v3n]QS!��Z�3|�g���+��p�6����:�l�;YCZ�������$/�DF�E[&��a�A�}�0�3!�n�r�a��$�9t�ʲ@Ph g9.�ۼ���%���vZ*�,�-�l��ڴm�t(�~�(1!g3�y�c(`7o�Gگ�5�P�v5<�1����w�_�NQl'�\!Ş���������|N䠙k�6՚�#�mF˱��9��qR��7�I���ʰ���R��xdq��Z��N�)2��]�W�,�������V��/�s��,5p���d�`����3:��8
��v�J���L@���I^��L�s[ZJ]���%)5�|�MP��cE��<��տ���p���>kذQ�>���S�1��o^�[kZ6�v�ˢ'�k��я�Oǉ��c�3�	P`m��c4�l
ǄM��[�V���Rg)�� �qu��RbS��\�A�u]�Z	���F'���ebf:� +*Ex���	"J/W 
�}�����+�=y��5ɳ�E�b�n0 ������q�	Q_Rŕ��^U˟fT�Y���1\���Ӗ�<Go
��-lܑo�t;nۧ0	 ��O°On�l��AF�m�bY0ICP��=[����d�t x���
��F�����L�V�HVD3	Y�ֱ�q��]�GRa{+���a�rV��]�tKM��¯h�:�C�I;{h再W鏉�s�@����6�A Z����إ>+�Ɗ֋�t���@�8B�R��N a���9���EB�x v�[U&�U�Xubs(��(��a�o=2��~�@yD�N]�������\7�>��9�ʞp�X�(3�T�f_��BC���x���=��i�p9M5��<2a�E��ۿ|̄"�����Ϊ�:c�<l��7\�J%�1n�r���o:_��{�Tu[R�-+*��b+�
l�
�a��K|a��h&�eIi�p%�ݤ����;�W��EYʀ�1�l�-�Ή�+�]
�<8�\%�f�F�t�#]���7�m��BJ�h6Y3����Q�m�F�M|���vg@��҂h�q{�6��DGX� ��N���/���NM�;��q�xU�*k�F�."$V� 1C�Q�}qI�eD/�Z�Ai+�*����Z�W����}��p�ɘ���:�̝�cX:Pjr�D���a�s�;�%(a.��^֭�)�y�,��:ћ�����qm����0z����:Y�Ci���o������H�w1*�ߛ��aC?��2SO� }{���Y��EcE-�,����reM{W������vx];�vO�-��W��F(#A�'M8�	J�5"���B�t��st�MQ
f����dX������Ȋ������Ү\W+�v�)��'U�� �n���E^bN?h9��he��U�i�+�m�b�sֵ���|�-:a��S��]"�M&�ǂ�����}w��V~bP{�[F�����e=i�uځ��F0&lթ�Ś[�|�ө�������>Rr�:�7����ځ-)��Ky�1��s�T�2|�V����;㠞�q�(+|�s�f��8[P�I'҉䓶��ڴ��(X,pq
�Ne�;��ne�7���ǋ+����,�4�K�<�z��#�t�Jr�[V�Z>e��]�G��L�2ю�4�M�˪���;����d���~�	\�R�lC�����r�yO4*�,u��� ���x:�A�~X����W�f2�|?�m.ƨ0Ox�(y��9oA�o|$A+ڊi,�FgYS˻���9��̌�Z�G��y|Q+����$)&ɘ�:�.`�Y���p�񪮭/Jͳ@b���K���*u)��42�	%������?}r��vD�΀�h#��Y*�Yq�/��J��2̫s��D�Z�8ـ7c�p�}� %%�I/W��U�>j
ғe��I�/�ؼ �,�F�g���p2���a���wR[���d�T��H�2�;��yܯX���P�b�m��*f٩^�������.��w���-�<�wy1j�"e9���	�lmt����_�ID��a^u�;�Cњ���}��<v���F{c]�򍽠d���a��Wa�q��y�WM2x�v���p�h,��!dmW�mc�wK�����swfH���mm��0BX���im������#��3�'�>ڠs��y�ͮZW%���q�^�n�E'D���	�_m��b�%�J�毉
n��o|\R8G��������E���}ؑÙ�F朻��JK���e�ǽ\��k+2O�j&�����;�Γ�	ۼe�6�v�}���L�ق�|`Ԑ�6�ڕI����7@��um�� �$��hM2.W�����T��=�� �c�Ѽ��x����%y˪eA���4���YA���a��7)�g��6C�s�K�	a�v�6�3���үd�]�`a���n
+�$����C�\�k����'BA$)N��0)��y����l�Z<x3�Ϊ뿔�jJ��~��oD
�/��'�$ʹVb���f	q{_��rM(���|2�rKV��[fV4�G:�2$@7n�[��؈�䗭�h�:�`�'	d�@��{~�>DU��J��\��Q�Sz�
�X�1��/���j�o������F��6\�ױO;vk!�(ޠ
�xf �*�lZ4�}� }Hn'�S��K֌�P�a��"��[�W�rW{�����q���U|�@q�:��($x
��������_��t���1�C�ߌ����8IGN5{ �����ƕ5������P��nrA�m�;�@�9#�(�����
�
O��01����D2.R�_�k�G��8�4Wx�vU�l#f���ŎÁ���*���,{|�uG���7?��Y�u��;۱�Y�9�\V&E���`�U�f�b�?�S\�ˀ5`��j�&yd���h�R�&�]�%�e�f�4GeW�Ε���#��cs�xP/T4-Y[�����.��_3�i��=�p@���������5f*;-�}z_��b�S^q��ߕz�bbT	(��KGl���>S�#��E��z�F׷y~��1{�0�9�����R��6�	<�%�q��`B�����Ut�GB�>r2M)���ѭ�M���1�nU�(,P]�K��8� :S����b6�?Nإ]�F��O�& +@�]C��=%{Z}d�ə0U"*b�Վ��XE����B���ո���b��h�p�5�p x.n�·�Dؐ�{�$�4��C��B�(��E!ӵC����{7�տQ~@@&[.HA�] (o�!>D}~�eU��3F
��;OjO���b�����)T��a5�u�����xL(���s(�1όJ�c�Z��Oܧ�0��!�;vm6��jЁBcL��hx�a�Jl~����+���u�RHG�U�)�C[Xx�?��&�
v�5�7[gmM������
^�5���b�=��JJB���nPg$�F�����/����1����RݰR�T�@���&��)o���W��{�p03�o������V9d@�	��gL��v����z��2U�Ul`��K ���b��{�R���i89.���Pu�c��zȃ���P��8iw���6o�h4�.k�����F}�̬\Q6���pM��� ������B�m<ia¶d�ņw�� y(�w�򉶈��K�Os��R��}
�7D�)��=�� ��"Bm��T�hC�8`�`ai�e0���.��@�`����`H £����@A7q�g���K��=��'Q�B?ZyEo�����\pZ� "nW�F�d��Gʂ��Xrf�m-�w������{k|����� �?^��`�K	� �v�ݱ8�0���y"�O �<N���%��T���*�`���r��㤽��A�̚�ש?�$�&"����):u������>�|�Uh���|�qLݐ���92�)B4"�i޾g�H��[��_�C���y�f'@ghI���4a@������b���J�[�VٽWF������1K)D�5"!0��������cV*|��������[k���E�wؑ��G򝥿w"��  ��M	��.�'g��645�u;>]����\�2v�6J7�f�����*��0ر�9� Ĕwe�gF�)�oi-�s3VT+���x�k���޴���=>7�U���r^jQ{6$*�R�Jٿ�(�K@�¢����`f�ӌ�Kn�������>�^в�
�i��"�qGʗx��\5aYDw�{3`~�uaӬkE@�m��|��n�����߮�\++�ߊ�Fi�����G��m�q�l�3�d�c`������a)����SD�-o�.�t�p1���K�ce1�b��	(�U���H�i���Hg���G��F��꒫	1�Kx��$�e�g���7Db5��9��m��Ų����6u:�k+����$NZ�Ĉu�L�:�	g�Y���t�����0���q��S#$-%}�����|�_y�N�cwI���&&�U���=�/wL�%�lΘ�4�ٜخUd���_+in��<>�G���9Y�ĵ��g+�8�WxZe���ࣣz�X:��,���X��TpYt�W/T�43��!Wk�Jh���$�)�<
���#�F���)��e�M\{�� {���F��s��*��&pJ�@�Ƕ=�ƶ��1�xIcS̈�]צI��R�u���&�b٩�׳�Bʠ[G���Sϊ�9i}ժ*\�	n�"��� �06ڶ��!�Hޣ��!�tQ%��I��Z�}h��M������zg����Y�G�n;���u0nU��s�^��T�[��[�����X����7Ϸ�)`��-��ONsZ� ߮FÆ���B��*n�Y�vY�Rj��&2;��^F��M&Е�s�ߞ/��#����h:{��b^�Ӏ#�V��Q����fBs���Ʃ+�#F[�=��L�P�G}�Y@��T7���%�?�wS�(%�:����IIj2��M���/