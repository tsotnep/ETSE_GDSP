XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+]-��7+v�愛r"\�b���=��+ƀ�wz'���=P�"v,O�^���$ҵh��Z��Z"��q��0	V��I�5U�n�i*��^_��u�3��&]��t2��cq�'o�f�˿CC�i�:��y|�C��ěb픜��
xP�;o*j�`��@ I��zrDOn�cy�
���D��OR����or2D'T�̆���řjIAzv��ұ��[o�t!k"�oE%�Iu�7t͊.3G���D�g��ݢkr�E����:�јΣ6��k�*����)Kf�@}Z� � �:A�X�d�L�+AX}��C�vmp12n�(��6������M��{-�P-8#�p�G��򒶣������P�.1���6�+Ly�9R![��]��zê�(n�_��0������Ht�:�7�	N�O]@�Cz�덲�$����
7e3n�:~n}R�t��!�#>���>
��\b�9�'.�����e<l����)n�
Y�L�g��.����h^\4����wlR0�Y��Of�˖��Aj֏�Ш���A�Hv��kv�	z�We�p��}�{O��6O`?"�`çNO��T�� :6�w�I��@�N�G�HZf��ܚ��I{��g�I�D��?kf��h0���3<g�u!��Q�s	7���d��o�r�m��ڣ}��C�������������E��xX��Ԝ����%Im�P�!��9�L�W6�%̉��� t��Xay�jk�>��dC�wm�	0��_�Xʺ�XlxVHYEB    aa31    1e40H�{�r�{��i�(����Ԃ�|�Ƶa#,�<2t?X�a[|6�i�}l�����F �����ъ�E){h�VC�[-�+uv�6<EV? �����R�جw�����{�����ȣ	������-��=�b�z n��~���)+�v�a_�.�(ോ�`��dX	�g�a��������y�R�S��l+��V�i? �t���^Q3���%vqzOR'�D�/��iD�������~Z@2��EZ�}ѵ��"��i�Ej��}&(���Gd?к�f
h��}�'W�$y-TN�S(z���k��(���3 z�͞;!���K&��Ӹ��bqf&��Ӕ�1�
��K���a9e�RZ5<o��<r�/)�/���q�ٻr��OB�J3):����;r��u5��3�a��	oe�4y!��П[D�*�v���׼F��#jvB�lB�p��\:�Uש�Ny|�;�A��c^�*�L��L�p��W?w_�����2��'M)�U�� 4ƆQ<=Φ�� ����/$`�=��q���>�d�	���P��]��
�b$r��k���$��蛊�٥���e�'���53�"����द/9�z&׶��t���S���(E�	� ����<��;SҜrq�ш��Y1�M�W7t�0h�?JR��+slf���0�X� �ߦy�(v����M�"I�<cQ�����th��S�cUS[�GK���=#�������	���5b�M>x̐��~��̍�׋*�8Q�Z5QB�B��x�<��
Pj�=���с�rsK��z��&P��Ƌ�,w�e�\�̬��]�Ɩ1eT�H�	����;�w=�Y��p�����W�,�g�"��{�e������
c��s��g�s�� �����(V��j\_�є�+0�<@�����J&s2���i~e�|'H�$а�
��d�59�,P^����{B��5��VG&Cm�E�6�::��1\���Ҭ���q�fÛ�F�f9�ӆ?��h��]�X}�e��ɘ��'\!��c��(L��ϲ���PHu��b�h�D��V�|��������z���¿�G܄��q��Bi�8H���*���?�C����A�N;ƢN� y����>x����F��2�+�j��<��| +�� ��jB������YH7�t�2i#�#&�O������C�B���7<��N�D��Sr{�/s��L�6[p�?���>Ia�Q��/R�F���`������XV`�t1m.S ��
ك���|�0ĝ2��P��vj��F�5�'}t��2���� o���� FD6�$�4-���$Z%ߦ3�)����Xa��
bre2f�UH��Kk���p����M0)�KE�DVk&���)!a�5�+hQQ(4�&Jg�"@F!������0i�uT���%��PA{��O+�>�wO��`al��;)��y~ޏ�I폌E�Z -=�RH� Y��Qe��[�����J��<�M�|:���5��O�1�(/�Y w{@.�gP���|:9)g���yfՅ���]� ߆�S�6Zn)Fp.�,��^�k;֣f�T�lu��u���[�_NV����3�0�tϵ��^��A����m�MDV\lx?�~Xf/W.�OF]��B��L�p�O	��˫w�B6� �ފ����U�Ȑ�b@n9��qu[Og�Mn��@#&PC9�U��2�	p#\w�Lw@Ya���7���v�O{_QJg�Gt�ز�)~p,�	׵8~��v|�t��@ɩ(1����d�=��e��E=v_,���2}F����K�X��4��m�I����E˭K%�a/��.����Cbj�	�hW!�f�?ď 2¸���e�iH�fF֗�D��{�vkE�v�lR0��~��|�1��)O�:3.O;��ښ�菂�շ�*y���%G�E��u���$)���b� 6o���#<��/n��@�x0t��<�z�Al	�T��2
� 0��#����7�k��5��o_u�f�	�؊A/���i�������0�2���C!�O���\t�~��f��w}^1��#��Ɓmc���$������Ln�D`sOVJJ~f��Y�2;��V�D��g:LIb4p>`G!w�d��E+wm�5��J�J��WG۲������v�͑��|�IN��c�h? �y�P�{�(�(1�k�q��&��F�T�7�z��4�Ԩ�3�v��� Smb�p�W���]��A�:��R~���k}���\� �(xp�C�`X�������=(�b�)mapLn-����q�-�=�S���N�`���}�� ����'2R�U&�NӡpճB�H�g�?��)!���������k�"��gߦ�x������U&m,re1�:�3%��0��n������U��ٍ�<]P�f2�:�_jor�Q]G��]!�)��w����,��m�DO���(���S>N�Z���=K<b���&c֌�� TCEe<��Xz@KΝk�iȴxmeQi���D{ı�|R��O���ŨR��#����'f�3+5���3�g��
 k󒋃�,Ϛ����|����9��n�)���q������yFdn����I�>z�����ڣ�P��yv�<ߕÖ�*c�!�bE��5��Ꮔ�V�2x���П�ɳ_���U%f�G�*:�4�2�t����G��-�I�[�c�q"Z���0Z�<�;td\�\��.g['�C�d��K�eb�Q���K���?n$�ǽ��F��/4ϱ/�F6߭E".�����=i��ΊkLrA/��ǩq&F'|?��w#�
 �\����� ��d\��&��́:zj�D�˴ l��B�LG��g�$*,����'���א	|�P �&���9�d�/Y�w&ڛH�2M�� �����W�|񂋽\�%9
DMژ��/����?�K}�j3��ΩU�yHN��/Y}�*�
��c��:hN��a�Lq�@���E��sF����=�!��36B��3#£�M�ߣ]�ԇ̡���a ��uҲDcO��%J����_�`�1�s�'�G��k�:��ׁ3m� v�(�xtpVT5U������M~�w�E�L��'�;����
�Ꝯ��=�!I�d��>D�O�d}%߳��KU�I���R��FW��h��]�pm����2OPe�G�4V|�֔�-ʗُ����1N��Oc#�Řc��Nv��������E~�5�_�Z��d���ػ���8G�ن\;o4�EN�e˝�� ��:��������x�J���>ʧ4xR(����K� �Mu �8>�`I��-Z�&�#9kT�h3���B!��¤������%K ��НL���bz�~ v�lՀ�Y'42|�#��d�����*IֲBh�&D�/�s�G ��m۠=T�>7_j��ܭ����_��neIȌ���:��ef��C�'�Al签h��t�'J&����k!����e��U�?����I�.�s-ӑ��Kx�C�Ę3�/=�^6��������1�4�%������420� :V���T��h�z������7�"���c��ٗ(�,J<�U�������Wh��a]x���!F�%m�LY�a]�ɉ~�.���mOY�dH�=t��`��d�C@����bJ�h�����gS��ͣ���qɆ�W��]3q�>	_y�`��Z}qd��]�����CTEi�/�y��˔��ІLX��g��p�θ�3�U�ߤ_��eʈ`Úހ�Υ���6t����ʩ�x�i���d}����<V����c�к�Cn�yU����u}z�q�O�S8�ۨE��0L2A-��T��V��J�^q`�$��v��O���S�5H����hS"DrO24.(�1�-屗� �2I/��ݻ{czqɒ�ҧ�)w�K����*��H<V���署�n�Ⱥ����3�*��y����e4�B�@ݲ�`׎01�IXTQT;��V�t]�gwXps��x��ۇ�^�ʙ���氏�7�z��J"��r�'�X:[t2���v��c���%�|~B��?d�?���;��_w4:Қ_�K��bwr���r������Ȼ��<_�Ć�)��q���
~)^x)/�5���.�jbCI�X��S��s�H�h���H��3��O�@�&ب��tm�2�!x��lktX��j��Ǐ�w�Q����#l����vi\����K����8N�c�+Ѯ,�P��B7��E\���M�vD��j	@S�)l����[���*t��HKZ�abA�˫$�7^�L�.��*�T�E!V���Y��5���ӽ����@�W�@8ml~d}O�2��MBΉ�fɥ$kIFѳ�)���ٰ�Q)��A�N2������X�{�3?���BIv�����jW��Qn�2�]|�َ0<F�P��1X�"�:�^���T!V����CB���i�u���.�\��(��׹r�&C�����;b��]�ȵ��?[i>ҁ��yH�����8ם�ᾉE(�PM�O�P�,7�`H�#���g�QEDi��%�$�U�0�mg��σu(`����@~ݩ�n9�A*q
��È�֌aQ�^SUn��7�.�{\0:}����	(����keov��Ka�2bS�(�*���U|'�逋���PΛ�O�3f'Ѓ��6Ě%M�}mE�o07z�P�?���-�lN6^%�e |��$Z6�Px�[<
���qc#�"F���n�@b�ԺH��4 9�"�Eo$(�n@��@ac�=hr��%�#;���R
�wI%�C��kӭ����q����,v�Fl��f�B������ ���Xូ�0P�'�a��}&�?*ܿ��+�/	bޛV:"��-�*;�;#Jp��-nU���vV��i�wBG����5�}�k�X	����	��m)#f��Dl��оx�U@U8[=�kH��%-/�t��p�dg��
h0ݙѕ��� �:����V�C���:����`�h�	/�|�x��N�['>��V��/�G5���"vK��|^�Ĺs�{�*��������i�k����2-���،t���k�Q^eb4����^��OsmCH�Xi���m���f�f���:����`�pVW�m�6����r�3�٪p��vBOQX�q�A(�.fa̗^�1Hӷ85���8��y��Ò�0ڹ��]t�F���<LK�-��ჹ�WQ1��*�_==h{�O�A�_:����짂3�z�d����^��c]��Bع�����N9<�1�wI�]�~>�B��O5=i��@�b���3�S�'g�G�k���e�������0Y*�b]
B���N�\m5+�&�
�.����x���zJO,\�25n���jī9Z`�}��p�IbeP�!�D>��T*�����
n
<T*�V��g��2�yyϧ�(d`�q�[�zt:�:P̉�x��|\�������و��px�6�:����6��ʙ'r���|�=�c��M�K� ��5G�-��\�^'2c-�Zč���>#As�����r�����}�ؿ�c�G�Sdr/˙���;�U2z�`_m,����35όR�j%2F����ء"�+���NXʁ�x8��z�px�0Jm-Ȋ�\�@�G2PcLO��]������AW4�z�z�������lǞ�-9`Y��<�)O/�9-��&���̌&�Si�X�	q{E�����}�?�c�<���ۈ��f�����[��0tFI������ w�:�-F��4�O���cް���(~ zF��P=.�?�˃��\���DXJ�R���
�6�S�� O����#8�:|]�lܞw��Z�` �t��Ǿ�[��FF��E=������}T�bV?ӽ�$�J�����o�ƺŗ.�����~	F�QrIo�Q���7��� ��;�	��L�Xn�%��8�Z�^��-�h��%�G3�ܺ�t� U,�i����yp�0�0�_�=J!z3ɭ�%/g�nHmE%+<<@QRz� qt�/�j�8�?!gH/�M�o	���v�In�ב𥮃n���So�A��r	-���둪:h�#>lr�:zPPK�FMDAj-h�����CӾ�Y`Nþ���Wnb&��j���;.��.Y�+oqC���X��bX��TˢÆ�Z����;Ի�N[_5�FJ����*:�=+���kc����1���h�U��\��������3�vK	��?u\]�i�@�rs[-\��On%��a�{��N� k@G�7�>J�A����n|��%2i��O-�32p�C�d8Ż���u���rI������uD���*]�"Ks�;��_~g��\^[0���.~��
����k�y"��S-p����,E��p$���(�<1�W�!��v���׬��t#����N���鶃��B2L{��X�)��aN�3x���?R���qg��dP{�i��L�ʽH#�A^�sQ�r�"�g�(��A���-[��͍��R�U�d
�h��C^!�ĩ3@���j%���Ʈ0���;�Ob��������uJ�WH�X�)��h��EyLX&�`�a�}�*:�mk��p�3? D;nx�����ʡK�\ݓXZ�t�$�Ҩ����F�Ϙcnd��go0��(5iI#�>�z���*h=�����ؼ��fb<~�0"@��,��Pm*3f0��A:L��#�D.5�d��=7����z�A5d��N�{�H�Օ�t�8�d|T2*��bA��*���^�B����'�5O%˨Ú [g��\��M����L�Z��`iY"��]�Ͳ�z�z��C�@�톡3V���3)�包���*\04�R�1�0��K�I~�,5�8'd��c
 ϋdɁ;o@+k�B���X-�ܽ��ۄg�O�>��g�?�j�FT���� $fb�����M�1�����h���<����}Lh���B:�q�e�b�CN��5��Q�4�\ċD�����?�870��[���]g�7NY�3H�ߍh#��ea�VQ�fli%���x�,+�x@�#~�.W2[.��D\��Kw�Ǧw�9���:���� g�b�f|�p��Čg�d����{�_�R
�E���O��F���`
.�X}ׯ�`׿\*�����^����c���7 �}�w�t�&ਅ�Q ��� @��$ĚT'���t
��&�~A%-����y���\ʐ"�VO��$�H�ui��_�f��x(jĞ	��[��U-c���Yƌ'�"���J��v����YQ1�<��< xb��!r��6#1�x��6f��Ik5\�ц��5�c�\���1>����V��|��K�̣`7�n��|`���C.����oy�������7���l��_U�6ԣ���Aƾ�5`c�T����c��5ێ�#�"�Ij��b`��./�����F�n�lL�"Ҳ0�$r�b]�qb7!V
@����S�� v�A�;ɗ��U�_̱UI�**6Q^�@w�Jw̎"�|���zGP �d�J%��e(�L��*��N��*-����Ix>�yu���H.DE�~�.a
�����y1�X�qj���4�)ܷ�=C�9�bf���%F?d��2.�p��&