XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8&.(+�U�j��_)��Y��7�W��nokQǌ��&eC�H߬���Dݺ#^���������O�����X�m���@��TTM���{���r#Q������ET���H�����3�X��#D��C�ZC����mp�!��7���gD��O&�~�����~�n��+�j���6�~-3�x�S1#3ϫ����z�=�b{#��/,u-��3*xL3g1�~55�X�@/�����6�fj^(�mt�/G@*g���Ħ�%����^gTH��� S6�@�CX��Q��w��f`�!�ka���\�U�l�����+R�c�������9�9���	!3���e�4�&V��g��bN�I�9A�v�-i�y��W�jQ���yLzT� �����K{<6K_)i��.A�@�>�(\Bl	$�v���Lǲ1��'�H#c!Qd�d��)�*����3 ���#��A�7�/�3������-����t�Ň�bc�d������ϵ�&�f쁳3ɭ�������~}�V<�v\+&.��R@H��ƛ�r���S%D����B_y��2a���R����y��+�a%؋����e�J�/O-W�O܋
��eu�#��R�ο�,i�LN#2�v�3|�; ���@!�6��0�ޠ��.i�z}D��Y�����1�����t�'���s�������2� �0�2q�P9w1�d�~��� 
�r���񟑞�G��I���3Ҋ�=�0+��`R��LK�u"��OXlxVHYEB    fa00    28c0.�gU>EO�9k;��԰��Ƴy Wiy����Λ�ͦ��g����X�x���������5n������xd�QVl/O���
��a��᧲�cs��,"]�-gl����k�г�Y��5y!kr���e��S��<�������}�[QVݞtX����*�)~� ��"��H�a�[>�����sz�1�*�ᣞ��{(
�"Uo������B� ��Qqd��YԲ�cѩS�
'�{�+�4��^M��V�)Bѣ�GL�Z�_�M��H�m�d�����/�O���ϦOL�#}?���G����b���h65�c�7�
-A�H�y�EF\Ԃ�]'��,Mi>&����k/9|L�Jj�vjE�&�Kbo9�0v��5!����ޑ��(�O�� �p�:��8�Zk�?p�oPZiO�"��1g�p%jz�1TY�c��[R�3�ܸ#%���xS�G����=�rS� ~±2S�u�ˬ8�Q��z��%d�����)��I"���朇1OL��ʍ������:%�]����c������Fs��Ķ)��%���Wр�t0d ��y_�R;k^��x�I��dh���E��B��#|.��F,z�j㇃�6%�Q⪂���!���;j��qBY�Z����/fk��O,���qД�����pQ���b��o�����L���q$0�M�S{N��w����g�����]qH�9���}�(��	�K"�r���V9
,'Dɍ�J4�����}2tV5��`c�l��z|a���0{aH�r)}Fmf�[���!�r�l����5��W���F��d0���b]�]�3Ь�H�.y��:���+����JqO��ߖ��[rt�~���L���_]��}�S�:�՛!�~e���_�M�E��"0(v��(.��l��47�?�1vI��3ܜ�;}ӿȴL�r:K�8�������c$#T����*�#~�j�X�Zվl�آ#c�L�'��hO
�C=����)' �,7�	���.��p�q�]�4O�g��4R�Ӄl�>�BN�!&��Lb�L)k{���ֿ�z-��� ٍ^I�`��d]B`'�WCf�C��\L�Ke�S��������z^�g1n6azy�)o��k1��Z^!�C�a�.��cf����G��;��㌗C��oV\�I�^��Z���8-�4���� �M��X�"��h����`g���1]�� ���O�=����i�Z�B���^	� &V���P0�6$�>јH�("45�3�Ǝ�h"Q�H�L-&��|R�Rv]fN{l��h�y�M���s}(ʝ�>�!��;ޅ�E�X19�)[�4
�O��<�t*�ӡ�*M��W*�6��&U։Tg��d�z�gRY�_���|ӻ��v|���j7��J@=���_�q�A�����7d���ws�	*w���SFLK�Eˎn���,�M��Q
f1�g7s���df|�7��I�
��2�r�z�������=
��H)y.�����)0T��"����k�P����S�_E^�ݝ�
��,�d+m��5ڡP��x��R���Y�qq�I�zPe"+�L����1C�Ѳ���Gr��������'��_�)!q�DX�E+��5`_&�Ĕ�0Z�'�>}�c��N���}rbnaz&[y3@��%6e�>�\h3جzf��ÚL���*��	p��>�Y��a���(e���$����9��[�:��������� I=�����S<��5���j�5M���dr3fzC>=����5���Zm��q�|jO��7l�Eٮ��QU�7~�0)�f�:�]1��0�c���ပ���:Y��p�9�$�	��0jN�+c�dfb�2�ig�}����+�ڬ�4
�4e�� 7.�h٠��<��hrp�R�ӕ�7W��_)	@�A@͞}�Z�� �y��8��%��<P��<����\C��T�U	��컌{G��|�.�5�6׋kYmaܢ��
�`q��J!r�J��9�a�QjBI^;{`1@%����(���{������|5Ǯѫ��s���a��T�`R�������:��Mm�9P�X���q��
>΍��IYK��}m��J[�������K�~]�-��	V[#<��-�_vd��Qq�5��8jwq}���ڤwj�桓���Opt%j7�X\�����[*2��}Qw�'�l��H�vs�-Ƒ+�����J)ƘZ��E�0��A�V!fz���O��ޛD�u�Ly;gO��*\x�Q��q��H�B�?�QZ�Y��F�b@}����V w+��J�u�=�Oi�#�v1��] ;X�� �/T�w\Q��|%��4���!x@ɥ.M����`�j�H&1���h�Bp9��CR{#�1
�z�(�?�\wH�j��۶my�Cc��;K)\K�*����AX+��E��'��lu
�S� ���*�-f�8,�
�=�yj�����:�5�I�z�o��ngh���0S��~@��e{I�i��@wN�WPR��Czf���KMDh�2}��٫�͈B�����`/��O ��!�����|�{���+d���^6����0m�n�2�"c�O��W�R��H�Y�4[PTD�UFTd�}p>w�xxg5�-��M���z��E��R.Uqݳ��ܦJ����~�����������Q�Q�5��x �,�����jԪ@��L3�5��֗������4E�� ")��:P�K;+J�3����W���W6Yv"6'�����޲�ʅGB{��Ѓ@#.�U���O����,�$�e����ut�m���(���Jr�?l4��>Rk�yLux��f����@�*�,�O��[��@>�IK�f���M3wgCT�q�9�❵����Z��t�`��}1޲��`p<�}*N��u�#2�Q�{<�0t*��8���J�/M�LA�n\�|L|Y��Ơ2��Mh;����<�Z��E��09+]�P�� �Hg��3�&�������4*_m,P��DJ;4[W��=����1���\U�?)�cW� ����"�`�=���-m��^������A<������ZY�h�`�qeEl:~�a�I�%�~�!�.-��w�(���In���-)���/����p�� �Q;�:31B�'5�9%6�Z��������(:���J���k�҃�H��.x�
�D���a�n���z��4�>�,"8�elVV�|��Zy^�*�`�oН�:���	��[5?I_��� q�\gyğ}�� �V䴜��!?ۡQ��*k�v�T�q�s�\)�:/Y�J��>bDteJ���]�r�I/����$5k(�o֠�	oFf`�XD"A��)B~8~aA�o�t	V�\�@K	ZeOZ�_#�7�|�i�Gf81o���w�?��^��_	Q�-0oc� +Rp8�q�nK�G�E�\�N'N��[��՛xa���_���\���)Q���lZ��N���u0�?��D��O�&��|�LȮ�Mg Ȫ��~2�h�X�����?M�9Z��A[�掟ft.U�S����1�y��m9pA��g҉0vG�֊'�y��������ΐ�Ţ�b3��xg����TB
�a��\��e`���/�C�W4a�~9�)�������+׻�Z���������W)m`��+ �������53}��j��y��u�	��o��L�w�9޹.i[*_���b~�9���f��E^8�j�=YY�}�Gڿ_w���E$Y����K��@�/��5�V�5P���E��(��y�++lf{Y����9������P����=�o�ߐ;q�
BYj�1�w?����$kR�(�s���!��WG��T9�����F����|j2����z��6IIdY?�SRA�c8�xl��l�E'O~H�����ß��<�gz�����:ظ�7��b���_yZc�k������Ö#��G@�R�ۧ�3V�7�V��=7����Wl��˧���|�?� ��
�)�a�']!�;8���c�1��0zm�c�ׂ7����yk{�c�̥��.L�>�T��u۪�SĠ�����i�����o��O���9+���T���t}�BG��V[�o\&hW�F��^" �g`�������!]s��m���V6��M�v�sPP�����t���:�X�� n�Z*K�ŕ7��Y\y.W�TU�.��Ɇ��>�����������q��Iu.��dmi�$�6R������?�Bq��Q5*�	l��D.Zm�d�����h=�ߎ�q�
�uI�^���C�*�y��̤���7�iK%�ں���@'x�_�7��ωڂ�`,���	F�K�p!p�dT��&���ڜ��O#ɱQ=9f�IT��p��&yť-P��ڃ����^��Oz�>x(U`�R~���I֨"�l86c���ĩz.x	��2rq�d��S�,��v������}|[�����0ұj�p��K��i�@��i�}L��� �����BC\Fn��CږPk}��q��c6(ˮ��2�XΫ�~��m2�8~�	�OO6=��B!�_D��Y����S'V�`v�2G殐�T��mJ5�U�8�����)�N�YE�N���D��k#1q�8�i�3;�@���`��S>�F���Pꃤ#7���Iy充��j�^�Fi�w�B��N��HYPǬ|i���d288�3X�nh�6S�6�w�&�_�8;E��ԷD���1����9M�+� �l9��O��T��QQp������B�%�h-X��F�Y?�Z���8�qc��}zs����Rbl��¬q�Z�SZH�~�P��-��"��0�_I1��9\��W#�g�кؘ�4I�h�D��@����s�����_A�:Z>>��_����M�ے��wV�"�hc����it�^����N	�m��R����JC.t��t2
[+�Of��CLf,�3!���gN2�h��>�)S{U�\mM��P:����W���*���k����Ƽ:.jc���q�fM�/o�x��F4��T
�w���Q&����gi��PN�N�f{����?�ld��˨��<d�j�:y�@d�!�\vê�'X|���+�S�9x����Z��/�<����%�>]���̋M<��쇣.w�%�P1��]��	k�#�[��$h�\-T;kd����J�إ-l��՗i���[s��{F(�LH���Rԓ����^�조T����I�5g{�2U���@���b�(�Y���a���k+�Rƽ��!dR�Ri�1fX�rcUݥ_�N�;�3�:+�d6�J�Ic���T�`�y =����ԛl�n�[eI�6��Ifțm_��]3�ٵ$��n�n�؍n�T���p�K���~+������=7To6�΅g�fix:�ש���<i�xK��mSD�1|Ar�2]�k�Q�D򣭂��a`�Us��0��Q�"pf�1҈|T�r�j���?��*�z\Ưv��̘��K�Փ ���RyYJ�u��S����A`��eCP����#�ѕ\��* ��&��}���AQ�{��v��=;{��6�s)�c�%fT\��Tq#�>D�/I�4�����.�� $yQ<;��MnT��@�γ
���&�n�D�@D{�[�@��n��8�%��2=P�ZJG�ڮPn٣�D	sS��ix��Y-�\g�Cg�F��m��N�Y�A�O/�ߎ1�����;'�ykǁd�A�qA{F��jא��eo�#E�{3p�xK��~���{qn���M928#��'?J���gp�ad�	��)�ί�O3���o2V�r�����1�y�vE�E���L=�T)�{����a:�K�2�iwhfd��\� �+���V�i�b|��
B�h�Uq�}��aK13��MQ=�{g�1�^c���&{�Ȁٕ� &em&~���5����I��1���Vdn�m_)���hK��}�x�a�֐^u�Ӎ����L׀�,jH]4��1�� ��6���Y儖�3F��g��y�`
��eĮ��^�Ơ |C��ש��c8��.+`;l��6 �*6���ߗ�j�P.�D�-'��^�'�V{���"]Ȉ4�:���h�Ӄ%?�w��%��ܟ�r���x���Ŏk���zn���r�z����*"�YY�=b�z�r���|�!Q��Y�
uX�N։0I�Z��ȟ��[�W����p%����^�R����щ��#�Z۲PP�w��jf_u�9ϰ�7�J TNxZ(�2�"k;q�M��jC�M��,�L�lOu?�6	����iE�'H
�;_��͘�ֺ�+��ym�K�AO&y�t_NKV�n�f~m�}-Dd����R�J��sW�۴' �)���ߝ�`�xӒ��ڍu���sD��4��Q2�Q����~ϪM����ȃ�/&[�d�9�3|yc�.`xK 8U�;�;<ΧA��^�Uʋ�?�	%�h0�騌�|�k�-ie�G��?� "� QLO��U�ԯ�����t���7F�q�U*/
�̼/�0���Ҽ�J�?�Yg%�#���d����B��H!��KSQS!!��nRP
�G�>r�C@�6BnV���v�-��"+%{�e����'Q��8��Mh�qv\�2��i:l��)Ռ��K'P������Xgj��Ux���#��i�d���p�6�5眿o����r/�)D�� ��q�\���R�n_�«����L����[/^�g�쑚��a��P�6|�qo�;����9J^U7 �pض��
��SQ0�VK��`H)W�������t�`�طᙳ�1��� �ZY[&mՄǂԼ9�Px bb�������q�����O��|�@���Dl�B���C@U㋿������ђ�!g�n�'K15:p>�o\�����`�&����G�A��`���y�q���=��#L뤯*�Ru�'�h���m+�F�~�c\�� �G>���#x��$���6Z��UIj���w�LJ���k�Oi�״6��Y����ݝ���s?$t�d��֗u	Ǫ�A`D�e��)A���R�����EW�����g0�m*V ���n6dw@��u�/����ή��6����d�I�� M!�L��P�9OFA�c��V@t�F��gq9�G�!_��t���J�"�M��Ո_S�w?�is��9'Z����I���\��M��>�7�tXMS�i=s�Y��B|��ex�28�̈́���]�+�M_��t�h�nk�R�d��P����</�UA-ݚ�	/Gjx,]M�	�\�[��Ci �$�W�����tj}H�f*���[n�ݺc���%��FVQjƉ�U�x�����'õC��W\R[*?ܬ���l�"�ʔjW%^�o��61'.T�#�]6�)���/]��ܾJ���lr)	%���+#|B�ܝ�A�9�5�$mӗ��j�u��)���/��n0f:PEq;��_PO{!h�-�}����Ċr�f*��3$ѥI!��zx��r����*$��s��s� ���ıSP٠Ρ6��l:���w:��ş Αi� ��m�=E�Z�/��pa><��6�N&#Ԡ�����T��Ҥ��{��E��3bQP��*9, U���"i��t.�h�� �9C�-�V0&8��f�ˬ 1��QLX�@.}�k�姴��?��/��
����d��"��n� ��zu?�n6�h���\��B���4c�њVFB�#���տ�*M��* ������k;\G%{(?X��N\BX���5B�:���\cՇE��e�a�<�ݕIУ��HpÎZXB�b��Ĥ0���W8�����<v���m;9&�]�|9%�X�Xp�5k�&*�]>���2�����<@�P����Ǜl2W�Yx�`��
�e~�*z�Q9����F� f�i�ʊ��d�r��mFW* ���;��<�ͦ�v�.PY,�h����*o/���yt�=C/�B����I�Q�N_�t�κ(�y�-!��>�M/���)X��Ĩ��9D��o��߽�DDՉ��s�{A=?��$LQ�� ��r,�	��i��E�3��!�A�)�Q�X�&W�b�D�}�Ҿ�,~���Æ]��.T���P�rdf�ib��Yp �����Ng��Qع?�`\������ę��P�i����Ru(�3h`����L*%�2��#��������9�����r��F�	��0f;���ⴥ����S�HD\"�h�_��Z�\^5�ǆ\U�:�	�3fAKL��lhPzaڞ�����y�B�����*��?ր̥4�~#���)GS���[=d��.wzs�7-���x�V���.1ȵ�so�C{�M0dg,���G�Z�:t}�zS|���Bb�8��ܐ���u��[� ��_/��Ҏ���GI?uOl튜���x�����?z,�nSmn�lP��v&�)́�6д[7����"`����^lH�UF C�]��\38�7�d���|-�Uޝ�����D�����������"�b��̝���i�'�o?}aC���SV{UJTp�g:��^;֠��(ai�u���f�ARw~������W!�XR�SO��
���>�)��i�Ia�c�g�%���5b�a[��9dm���j���u)߬�^�3����E��o�R�:8�[����*��N;�	E�#�tV�=�9��/*�.LP��.�,ɮ#���PN�����	��%����#��M$��)*����m�Й�@!N5� ��$Qr<^1��G.��@h����'��Q��!vwW�Y�UK_0S�7w�t�deW1��\���Cʼ��b���*�#�N�M\h�Ţ�ϛ@�d4XL}�g;��6�� �'�;�����"�o,bZW�{?�;N�"�*v5U1?��iR����C�y(�tٺ���O9����vu6ñ�<�>�+�V�dh_C׈��	���(��y��F��9�]#�#~t�J�7!$�I���Hύ���F�b���᷾Қ���@Q�^��N1�||��,R� ��\P��
��6�\�\�"�9���8�qW��>�T������K�)v�,���#��Y��������WX��}:�'|�P/��� E�cw(谚�}ý��l����}p�(?3��"ꓗ`f�ʼ��������[�	�O���}bƀls��r����}pn��#��T'���xM*���{I^>�=���
�j��ե�O����Y~��"�A_m3.�u?��p|�"�ݽߧ�r0�A���O9!�� ~��{�x��l΋�oC�����cC}I��{P�S��Z���jּS�
-��Q�?�ֿ�^����ve���_�et�Ae@�����,�����DE����C]ލӏ�p���9� ��)$r�I�x��9�_D��1-@aO���(�(�)Ĩ�k�G��}=��˅~�,�������R!s�g������@�L��䘸�[!�J�Z�)����H�1�U7W'uAQ�Y�`����΅a�9D֔"��,���;���K��O���G*ǁ���W���O��!g4S�V�u�'��otFWkӆ,���U��z�����]%I&�[��3�m�S�a}�6�zB(^_�[
S��=&)I����~�碽�J[U�y�T+�V����	O ���"5fY�q|g&t�k��cl�354:Y�!�k����tS��2�{x]���s�dW-���B�cP�+d
��7 \�2?�)�V��+���*�e���q�Wz�(���������sB�)��z�A!*���^�6a�w���͉h��ڿQq�d;�0{c}C�m�E(sm��:ll��X�5�p�ኅ���Kw������k�GM�y<�-<��01+��N&q�-��@��"ǐ0�͇o�4i�����3Y�u.��>�s��v�(dx����_��ʱ-Wi�{,C��ϵ{��m�2b�K��3�^<Ng�������b��ՋOџ�Hs�i�ҵ��"�=ܪ��鋳G��&��:��:F�ގ�����=�G����ߪ~�i�s�)~��<�π���o��ߤ���|'���0�*j�
:1/w'�dgo_԰��rlW�JB�t�7�FX���cd	+���1Ru���FUy��>'`�*����p�$��'k�ܴ}�v�������l�j����
ƃF	F�XlxVHYEB     896     280-���U��X��w�j�(\V�a�א7��_�d��I<�:����[���lc�p����Q�\B��[:]�
��
�Mw�F��p��c>�\�S�����%��8����5q&�;؏��h��lW:r�<��Pe��'�Zq�0�O��	��ݭ���<�U�YQ�yS�R=[|�\�;C]����P:�K��V�c`�x}�Z�g! ��͚��jߝ��㥵�aZ��ncw}8�{��!B�
7bB�vU!��ỸHV��*a�T퉇��I8U�`�S�Q�nh��us�[^7�6��h�н��e�TՕv���w _�W5��s����P*b=�ۧ5<�w�K����u-����T�6V��V�{�# �2{�O=n����n���A����S5�"Ym�x�U�|p; x &3(��"�PB3=5ݶ.�W����z򓌌������.�繴�KE�?����������j�쬟U}���Ŭg�˙�kop��;�B6���ЕE)�U8v�.F��o~�yL�t@%����&\VcE����x�~�O��Rd�Φ9���8Zpy3�l&�xJy��Q�c1Y5_�?��I$x�r���Z㈤�7�{��0Ou��.3�3U�A|šR�)�i�.���