XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ۂ�l'(k�AA���������rl�t:�ߋR;��_��|*+�^��A���9DF&{d�����Y'�T�:�aX�g�Hg�6��O´
��ܫּ�ja|X�L��wt	��v��4������� D��
���n�{Ļ�$т�v���^�uu�.�-��m�ۨf:���F�;�*���\�s�t���@H��ρ��E�M�hk�ŀ+����#w�+���9�g�/�©��U��l&5�laM"���
&���w�;������ص��X�����:���h�%��f�n�<P��8�i��כ�Y�����s���1;�g	�M_�k̙����R�CE�K��$����,YF@Dh��|��S�L$_+��
J�*��K\^��!��"�t��U�t֣=����܆��hI��~��p��p=����oN�)�*��J5�2�(M�b1*��µ�Bgf�7�#d �=2ɢF��yyw�^��Ð���Z䃇��"��X�p�h*qU�=�20����7��,��G�@<�[d��-�:u��#� ��	v�`�-q�ȇ������8DCBtS�)%E�S�\�8���:i�X���G!��2�Β�rQ�8P�22L{�,cZK;_O`X����+�	Ҵ�Jv��F1�#����c�q�z:���]�y��wRT&8��*e��H�f���c˲֩�.�����9IR��G���+93`��Nu�-qə�	�Cg�(HG���"F�p�W�xRw֌XlxVHYEB    fa00    2260��j\ɴa��N't�6��T���Tv�)H�PHm[c�"	đ'���i�.D��̴�Bd�G �Gd���&T"�S�N�--�����O���il2J�+,)в���e!xwG���#̆�Y\��t�Q�$��;�PL��]!�(��q`4�o��j��"���?�Y`2I�@kjg##��0D�_(�:l�e��<�fR&�á�~ˋ�j��*���,�#���ۄ���ٮ�B{+���PC@7�@`r���٫��_��������Y�5nh�"ݑL��7�eB�N(<����96��M����3p�/���"�N׵#RW3����6�q��+��f��{�g�w��ݸG��l[�: 5�}�9�4��]�H\��\�[���2˓�|B���?VZ~9�d��˗�%yq=+�Y�"q����4-���Ӽ�����h����Д=�շ��j@�#�I�ќ� �?�r*lXHd�$�:$ʏ0�QS�����'Q�爠�F\�6�m�Z�2=@�vf?(����xzF4�|����������r!��5���<怪��.h��V0i��&jq܍����xq��Ӈ�6��NTC�h���Au��J��H�gD��%���buW����@���D�j�O]`y�8�SH
]r�]�IT6�i��m���0�[)�f��]�.b�+s�W�0t��Y.̧ھ;��I���+ۑ�.�}�01�]!�����H���qzN�>�à-u�n��^A�/�@��M�q�G����f���`�c�Cg8�PX8e�䟖�ALܶO����TO�I��]$�v���('����-�Ԗ*�3Lo��u�纨�#���<���Ӭ�O�z�'y��l�Kq���pۏN�"p�D�-�B��ң�b��ngC���9�uy`��?~ԣ:���5��P��۠�t�	o��}9��P�-F��|�2�XMڄI��v�ㆭ��*��`O1���:·g��;���0����d���S_� ��v2㜜,l�5�z]"ZbTp3�����8�����*D�&��\a���4Ùl������;NR�M���k	�
��[$2�l��NՖ�K?D��m+4�y�28p}��E���; d�4�P�������'NL���� �C�l9����*7PJ�rj�!n�困�P����cͽ�h&�	-�e[!��Rn��³����{�0¥(S�m��yr���?|%ԟa�y�r�W내'��ۍ�W�.#{<�Y�Ȧߌ�}�P*�B��d�il���f�ߺ�VM�6��i]0/B��G���=���=Y�ڕ�>��Y��ďbČ+m��~�F$��v�ߙ����u�{���e�e�$�z/����p�>E���j5���T�|OyJ5m����]�;��Ps�m [��@�|e�B��{B0/��W��Հk��RW��&�\�O'�!c�oΕG?�`#�A����D�qQ-��+�O��|/0>�E{U��==���ĳȾ{�A�L����I	�u��5�9�&��֧�%�X*����f�ۖ�2po�����蝿�z����TUȝ"�{{@��$�U����Ƭʇ��}�a�ߟ�">-ZO��əC�``sh��{��J��9!�	I'xF�����`ɒ[m���D�����q�o*B��@hl{���oJ�˯UR�7{fGJ�6@{�����ӌZiY=�7�����I-k���l1�r�U)�a7���W�@ر����it��p1��
#A$� �?J$�Z>�qh�Z_f�y��r	A�2��r��E1�P���+(5��tL�9
�%N��-{������m�T��E�P��(�E.�Ҥ3��cO�X^�
/�q%ߍ÷R󝔇O���p �z�hh�1�P��vY�C��5�9�t7a:C5�,��e��B���W��`f�=�M�!3d�(y��(è�imG�!�������4��F�����li:���P�з6��	6�(��\�~YE�V����n^7�����i7�EG��I���X�K���k���T�����l-F4H>Tc��ڋ�7���颔��\X���3�w���k�Q�#r�}��{�ҕs�"��&�ak8|��%5Ɲ{ �t�� I� �����bq�d�d���`q9�r�1?�K�����o�rB�}@��ZMqV�8����O��חE瞌2ҋ��f��/0'<���5^h=�z�b�-�˸7y��pK�����<?J��:{NSu�OQ9N	s;f�YS���P�m�q���(��I��j��y���3tT����3��`�wa���$��f��[��Ø��\F���۠�ݙ����I����riT�~ ݥ��)JVy��,t�����p�۱&�E6WLlt��V|�1�
#/�����ۂ�p�-8�G5D�sv�yŷ_V�w���
�5�f��vG%0w���-�?�kHM�������[ٛj%9G�E��m$�[�"�)Ȕ��Y��$�;���(2��P��I&�2&j�W�_,Rb�'�WZ���p[C	��e��Q�aQ<+�
RNe�x�$�t	{��I�L��Ӛ���� �@7M,�����j�>�����R8u��nFtع��Kd��f+�ʤ�f@Y��]@?��m>�J��;P*j���ʻpɫ�]s�r藘�Eks[4��=6 S�YOS[ͥ=��$r�B�.p�? ��m<�pؚ$�c�dz^�!+�����;W�%i�Ͼ�W�]�4�.UV����к�s�Vԉ�B\��r��/�7�Ϛ�w�&9M��Kv�Q(��R	�~.��Ģ��Ƥ����LN�O)���m�:Z1ܝ}�h7�`�}��ģp���^2��=<`��:9�����5����%�Ƹ����;`}]�hKB��v��$\o�?���
ƳqA,��ZBZY�Fyo�]I=�4��j�.<~�����נ��H�){y��7x��Kt��Gzo�� ���"] c*s�u����yFF�W�I��Qɻ@.}Ņ �=��~FUw-�^�p�mDI\\�f��O�~DP�z���i��+�ƈ�ep
c4[���(��� ��繴�}���YXmAg��&�A|��K��+9l�����\��"���`q�$P/���N�;�5��[�o��b�+�w?��q/>�����s��Q�(�2��,o��'a%dzI�N�����D�{of}�QmP~����}��lw�ud�h��@�_�wb.������F8�����N���I��"��z�b��R���	I�G�(�Ly.>�a0��N�YL;Q��$��Lk��x�G��t��}>�=F*�iL˭x�X#�j$���l�d�V�,��<����.5�q��T�ʶ����A���zԍT>k_�ҡ8׌�u6
b��Z�G�T^�}�g*�jz��ńw�Fs����ſ��5c�['`�ɇ��f��M��
FΏ�z}��aj���"´s��1�5昧�rdë}�F2뉪Ӏ,I\HE���ǖw 
�*��a)ys7� '��å��Xܸ�[�<Y�'�آ�}.OO.>��	Vs�(�@�[�a�Ĵ�^�HWYR����5�Z󿉗pH�V<wҖ� ���6<o��1:���+���m�^�I�jH�7]S8u����|���+�F�o���ٙ�k�yǗd�Ζ��t�V���?*ڷ��	ˎ	)�۾�u�,s���<Wܓe�}�x&%Gxt'U�o��Pކ ��lGR�I�nuc[p)���*�O��C4�z�ڙ����{;���ZS��)�0���Rklz\^���꛲�*JPRv��d/v�n�@+b�S�Y�Qa�x\�i��	ל@�H��n9:��Y$R��NR�WIr�'�"O��Tv�<�ûe��Fŝ�Z��O�^��o�Vǵt�5p
@-r������|�K�x��W�(���������;٦�v�w��n��-ʼ�E���� �լ���:��I�>3��x���D��5�Q����0�X��j)]%-�o�\��k��E���ro��E�0����j(�uʍ��{=_���3�-f�{3KZ�X��ʴ����E䵨wv!��8�/k���NFw~w����ؘj.ʳ��U��9Ϳ ���|���� jܗ����P��kf�z�=q�~���^��I�N�R�+Wa�}�8Yc��^�N�͕�Z�F-���a�<>�P"���+���jo�H�QI+'s�w�(b-�m1_ƒ��i��p�w�L 3���(���-���K���*9�1�$LMU�@�虪�M�Y֋�}���oA��DT8!�CB�G��!QP���5k��,0��H]'�sn�9�1��/�+[9eW��|n�P0802(�	�α�Gީ�%X=�B�<�� ���!���h�Ǿ��'���֕<X��>G��:X�v��)E(�ԋ�E��5o����z���ngsmD���uD���pw7�������D�3�㐟�l����N�V;���5s���7�6��;�����ON��n�=�W�N�??m��n����U����U���/�i��;�	|չqL�E�XT�e��ۇq��$�|E<�
�D�W�ϰ�y���S�<��_&p�e���]��/v�\��z�-����W����N0|*�͠'���q�Q�^���=��q>gr	�Wy��]��f�!���_�UC?Wej���א�#bo�:�I�k8�דZ-d�W��\f����;��<o�zHH]l�`�強�\NV��u,�DGu����h��Tq���L��)���M���
�V��r��+���a_��_�����Q�m��g#�r�]��y�`���в�;'vN�
%=-{x�h U��2��l��dY������bQ����[��n��x)����(���;{re;];R�v0���io��F���N�x~t��?�W���l>N�[�O���u��"N]9���?ʔ"�&�� �'�٧�KB��`���j��i��q�+��gי�^X!W������g%(�4ǍMFԠw�K��$�z�g?�!KП)�[��%�qM�[��mbyl�(�wZ�Vo�f�h>��n8�OF����侱a�v�%5=I_��yQ�P�IN]��!#B�~��N0�b �b�b0�fS�L�ʑ��3�ܥߩK�J���PH��Y�w�Ϋ+�+;ό���+ 1��	Ͷ ��@z���v0)��̍�Hƴ�U��Ւ�+(&tk���΀<7�]��+��NO����i�U8���Y����J��@�Rtd_�� _Z����Np#>��L)5�MCk�X�G�F�Zl�t�����Fy��W�#Q9;�P�|�h�A���B"�F�W"?'e�����y�:��\� t�=���y�/�l���+}Y3e��m���~�<�{re��NV�&�e����G^�-��z�*��n��:j-��p�c=�o��a�r������e C�t�a��IXڶ���*��~���϶-�v"�8щ�el�}��?�"���E���uމ����w�ld��x� m;zX�bV�8r�4q�5?� �o�MI�:KEp�_�ʘ�0Pv\���na�O;����#�d)2XiX�8%������K�+|���k�\�\�F��M6d��}<��m6��9R��3㱁ќ,�2���sZ"��v5����Q��X2*	!�)"��y��`$y�0&n��;E>�L������(J�['K�W�m~�*>�H�}l��N������BK��o���
m���A��%�'OMm�a���U�"d��V�wKY'w�5A�SG*�~��ou�	�CS�p�v�l�����4i@)����a¹�|�4M���I&�In�V�]��;\��`��'a1�~������.����X�d���j���9��1n��ˏ�f?�N�%���V�4���O�v�u�wm��m�
�"��c���IM�)�i�/�Q.0�AR܁ Nc��/�h����ߊ�0c�&\aS��؞�f����A���l)ȫŪu7&'x�%B�g}�Ġ��%m
e���ˌ����H"�[q(Y[��W�u�~�?�%S� �\CD�YA�@���{1�>�̆S4��C$[˭���\8��n;�^`�dwK���CJ�Z)�nz�!o{
C?}�nJr�O�ŭ�Ʀ��|S�'�2�����n���2��3�R\�CV��N��E��=��1h����ߝi���چ��'�!�+@I��4��(��Ҙ�cBo�^�4��c�D�,<�S@B�ۻ��*Sc�A}�+B��x�0p|p2��_�o΁�*�n��z K���Ug���hx�8A~��sf�صhп=
� ɏ(A�p�lkz�0v�iM�J-Pݙ
�j#Uye���ݥ����x����GrO�$�ޓ
��l)�N�1���� ��/�P:�I��{\Wf4�ld�.:��m*I�I���$�-j8~�:�UtY|*`�O;�:@�dy�2 �ȡ��@�TEi�o�:�U�"�:��u����F�^�
�nO�Ӥֺ��Wuʝ
Ns,���n���,��zV�R�K�>����i���Q_�kiyA�z��S�rh=��k�I��[�jS�?��/��|��������5�\��&����
F#��$�AxMn���@c���c�6��[]�n&�qB3:���,/����vƤ�>���0%:?ӈ���{8d�؋�['Zԇ��G����j��9��S{r_����Ԟq�I�&�7�#�
��R���H�>�%_��f&��Zl�gfx�(<�1�j�<Ҕn�f��
@ }i������C�mh�z	���k����@u �n�P��ZN��bI�7j���pJMQa��)�����|�ۂ[_`jq�3��&���
<�Vƙ�&�~�}y����*Fe��#�I���wA���/�:/@(,���F�?�G]gW������Q��g�fG�i�j�F|��*l��0 �PP�\���0��po���)thѷ!W3��Ɯ�>���f�|~��͜gH����Ђoӆ��Ş</1م�3syl,��)����0%�oB�pj#���+�AQ,�n�����ҋB��\��5��.��1\�O�+/Mf��N�\,���R ۳u@�&y�^��@��,^Ba�Z��׺�����յ�-$�|!���4���l�Bo�P?�j���̏��6���.�n��0�n^tos�
��o��G�Z���,���?�v�Ƅ��t%k'�nqZ�I�����rv���HNav��P�ڥٵ �D�/|��'x)�R����-��1��Un��=��9�N�[��/ᰩ��D@�����^n��{����R�h�Ci�ډ���ȡ��r�3�&àp��h�!d�p7���*�9H '�:��%��T����]j�����n��T�ښmX�q��D��;�1μ�`��~i(oe+��L �/�~E�9����Ɩ�|矲y+P�x!A�E��֩y 5I�ݓ�g�>�$یg���Н����}�!��zx]�4����mܣM����ɤ�i^�#��!FJ2�r�Q�z�Y�����\���=�	��� X2`����PWJH7.e�1���+TM�dJJ�ohT"�rF�r�U�1�3�S�+% ��$
Q����;�̜Xݷ�#e���୚���՚q�o�A�Gf�@n�L��o��+6�URp܁bV���H�\��᠏��7���0�|�^/��q���bxh��=#U����␞_��U��n�ח�z�oM6�x^Iˠ���c!��g
��T���)��8]��t�>����Uu���/&���;p�#L4'���T �� ��G�[d��,]�譀e
��
nȍ3� �%�w�5x��| �iW��rua�a�xq7�DC������: ͮJ[��;�ϛ���`pY�18�cF���r\����b*Y�G�y��f�	�̋
&���5/�0wN�ۚ/0��⢣���oFo�i�n�a	�K�L�n���_�ml�����EB����x�%L%��s!]�0�-���a��t�È�U�7 ��[�wbzu��}��{GHD$��]�*�_�y�>�U�p^ %jyY���w�Y���A�[����v϶�+��(��?�]t֪Cu���grO��sk�Ԇ%�åД�H�B��YM�l�C}��6���*�%�41�u���I6-��F�ؗЪ����vW2Hb��9a��/�1Ҭ���(��^qF�z1�� ��6��3�i��a �d��y�P�j<�&��u��tI��,�gKj�4SD�YM�Á��U�����n��-L��y�&S�{����g�7V�P�T�,����܈�����F��Q�|�
�7�h�Fr��q_].�ҥ��/Z�y�`t�c�k��[Y�`<���(���,���Bw)��2����'���|f­S�OSz�=�=MbP��>>���ɵ��=�����6n��I���1���уa)�*ܴp�۬�(Vi�<%�A�,Ǟ�|9���[�o��ゕ#���`� ?���zZzO��g� �0�A�ߥ�|D������OuƧ�V�4S�bL�Ehh�)j ��!�
�`f�
o��_�<��=�i���'��XlxVHYEB    674c     5c0\��Ѵ`YI�l�Cȼ�"����m���L
� ���o@�a��W���{8R'|��)�W���ݱ�d�
�h����33�$�[Y,��� �G���&Q��$o����t^/^V�6C6̛���˖�%�����@�~�b��#�0(���ӭ\] ҏ@�Z��ý��~Ƕ�.m`�Y�#l�ȵn~�\q��խj���ٺ�A��c@N�N)8����g�i�Y+���	=c���~�#��k'�Q���y�?7f��A/�cRW��C���Ji�V?��-KjJ�h=,�̝b3	�����rr0`$yz�j���}�Es%�m� ȱ�۹$9���������KxH"S���R�4#�s'��������9[QO���l�m��{�֜)�D����{D�S4zҥ����+=z@���q��?&I��A���-t�{g��r��zo���aԓ0��r�AՉ)���B��f5�E��n�KE��l��gi�(t����rTr͆t'�LѪa$ F:xe̿�6�W�B�&Z�S���xQOxf^w�(��I@��5-��(wX�'�Wj-�W]��5����\��R���y��!2x�4�;�ڸ��]^��N�1t>	F۟�^�9Ҧ��)�]�yZ��8�����|��5�e�m2�D�Z�̿�`*�9�權�V�� "9�	��9��:Ic��I�����3 �叝g��%��)H��W2�[���+�%̧�Ŕ�Po.m�5��j���i�UH�"��̎߱+�ByWإc�?�ݵ�A)j�v̓��(v����У�vz�1�:��.����8�&�>k�����6(�/��7V;Ktl���kKx��g*L��x�q���5	�#�w(��>u@bu�2J�ű��ۨ�٬�rg0�ɬ+���k��~�1�~�G�ۑ�� �ew��,�y͢�y�+�~1�ِ��+�����Ah�ּ���kO�Z�|�V��U�!��0�>ɎWxm�T��c�/�1�r
g$�r��L:����B��f�Y���TP�0�C&�W����-��eY��-rטԆ����_�|?��,��x����ط�j���xo����6^+tQ�DN��ْK�'��'�;�

g�E�eW���Sq�R8'�F?�,�&&�1jè/��X�ݥ������ay[��U��I͇L���Ӊ곹HYJ��K�TpE�X� ���AK��H@��qS��ʄ`u�To��(������[�����{i��uY���>B��%���m-�,�	���jFꝨ(aN���I�s��Ln&a�a]���$�h|����-������uܾ�\�a�2�wC���"��A������l&ג�y�<�Q�s��}W�D�o�M'���7�ǠY%y�ߛ��@�f�qU����iz�3��I5�z阊��������%�Z&zw�,i-����$�d�k