XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^!U��Q�_����+��� e|-J�HH�}�͢gUi�x"��(��7i��@��x�;����jH��[�{c�	������&	�px�՚��0添��T��TՈ�Y�EXlߌR���Ӂ���N��OY4>�_2�`�ڎT�X�b�u-�|��AEx�������Bz�R٨�"����1㛭��Y�P/��l�*������Yc�{i�5�h�2���d�}@c�)����*O��L�Z7���P���2a����̢7
�[�\�pZ8�4d�%����E��E���ϗx�>�VRg0Nd���>¤���+1b�#l�a�ШM�M@8{��ZG~.��&3�~D7Q�?�}�P�A#c���}�f]@���<��c�Q�G4���P�P�7��@s3��3��sY؞ӝϬrH+� }�P>hb�v������5��H��j�Y��B��}�$IE�>z�a��p,���\��.��
��Ji*���z�4nBa�SG�ўCy��(9�W�cER&IQ0[�E::�� Nb+�a�B���1�&캸�T��d�.�m�Z�l�r��F���N`z'�,L��RL˲&�kiU넼��p�q;nV�{���ͷ�}�Ȟ�v|[�V��Ǟ��!��(ݴMWI��WWPQ�k��ۨ`��b���[�^rAW�(�v�/}���Q-��Ј�J�	��<�����=���⇮��j.چ�}��h��ϻfQv=_}��n9�S��2@t��5ھ��E�4���Ӱ!��}�XlxVHYEB    fa00    2480��[0���%�.`6(�z��Bu�QU�8��������I����@�`k�ѷ��,K!��� ]W�����	���!��G�(E�)sZ�~����G��7�iŒƻ4����q�j&b�1�[Z�|L�eI��W.a�s�\�l�$&-�5P��+�G�����M�P�1�F9Ю�dz1���y�pGC`�Rm����6��?�}{�<���	#U���!�G1���J�� ���B\���X�R�}W,י5݊$0p��&3��9�E��ە5[J���=�Ӫ�>�5W"�1"fv"���A��t<���h#+{#��w��Z"�2�������G��[0�2�P���X�u f,�v�%x`l�I��~;]	\�fp �?�Wz���~��"�KQ詯��dqm���2ȴ@��;�:F{OЍn.a~��.��a9}7��N�d���>����;|N~K9��-
����n3Ez`N��	�o��O�6�p���"<[ص`���m�#{�.�v͸�h"�0�Sl#��q��"[SeF-�����M��.
����l�v�d�7)!���2������ŷ>��`�X���?(?o�����ߞ�S[�)��r�2�N5�mV������@����7�H�Fw��:�m&K��M�ܶ9WP�{xQ�q�L�vC�įv��g�;�tb�`�Ug�~Α�?Pܡ��R�2��5rbRc�?����U ��g��iՓ��p4������`��g�jk��04;�WƓ�3|��'>�WZ�G��gF,���^�݄�>'��D���O)���u��
���>i(q�p���H:7*�k\�7��4{���q��a'����;J����,1a>o���Iq�Z�4��-�!X$@�
���=V��z��S�X�3{��I��z��i����8�UwQv���Y��1!;8��|�!����'����+lsÎ_��iN0��-'H���¢�Fkh�'���9�'���0���A�QH��{��vx�4�.����kk~Yk�Q�>�(�U��PZy��	 a�T7z�۴ss&��Te2��H�c�=[]<����<�Yq�G�\}�_
�t��<j:��?ب+���R����f��}/_@�sM@�@��c�~��WJ�j;�<����Ws�u��n��O!5��a�ej _`�XI�%���{�=������4Mϓ��6��'c\�c����������3���Q���%st�m?HR������<����ס����	鼆�a%��8�ݼ@p		��!{���Jc͵�,������ϱ����2'�Y"����%,�ھ�??=����0B�?M��<����5 �v2R�N�<��~"���K��ʇ�yW��m0��A�0x?��}sI�W�=�Bj��@�*~���渔�p����ߢ����֨$3�Uի�R��E�bg�Ӫ�����?���g_�W��։�����p���$��rH�n�@;��X:�=AF	��{���Ȝ.����n`��Ą���N؉C�;7���0��-����N�/�Z�p��7�o����~��v�**�d� ��ό6�e�̋�B!��E��Q ow���͹Gt]^�h\ß%���g����bެ�a
z-~��H̶���tr5|{+��w��,��KL��5&��*tt�hq�]�7A�t���Xҫ)&�����fD��CT��6���~��	r?���,^�8>�b�X���n{�rD߳�t^9��[ػ�d��2M�:��ʒ��D���8�橳/#�v~a{E�թ>0�0к�+�«o\�x7�n���gs膤����c��{¡��~��oP$�bFQ'7V�3�^o쥱�~`�+2�?[����(%������L*�{C��Q(����\�~��ɍg)uؽf��ȫ�E)Jc��	'lO߸�o��fo��t2��=9�� $�вgٔ�%�>�~�u�ӏ������hW�T7�{��D?�d]��#��s�B���;�HA� r�k�]\{�Ԣ���V!����L
?�K[�X;�(�+M�k��#8I�;��M�G�=y�Q�A��E��̓�ݽ��-J��wlӖ��X��;e�Ѫ�K�pD]��
���{f����{XK!�8{_��;2�Gl�2dt�36�7���]�~ϯ!ѡ6\P�W�>֯�..��<��sv;���=w���v��Y1l�����#~�п���_��0�(&�J#V4�?��.}��ILn�N"�,���s�λ�o���'�{�2���6�Pk�H��crl��aQ��cx�����l��s�/kT?����5�GMZTx����f��;�񱕶H�V��KϩY`��{�Մ�q(�-��G�ڦ��& ��s�P|^�� �Ow3V��ZX��k}���b��}G9*\_�gY��{E�z./R�_#��F���zn�ْ��`�Y��uS)F��

	
��S(�F;�����|��j`�!g����/���͑��Ǉ~�	�[ �̜~�n �G��g����J�(���J"A|@/�G��t��Ǌ��}.@s�Ɨ�2����S~�ø�M����W�Ѧ� ӊ��l���7������z��	��ܔ�N�	s��_���2�.�<�J��>��Y!�9�{���[�z�����	Dh�e|�M�&h�U��շ��$�))����每2�\b�]v�o�AV��G�Ny��̉����\��ԕVJ:��֕�[�Q����|�����\ ��9C���<
#���T4ާ�&	e��>{] �g��a��x��g�e(��_c�X�Xp�r��`͏�����G,��$2I����'�4�O'�Z���xF;�J��[��m�o&+�2g�Q�G;)��R�B5�|��?�b��*ἇ��h�C��|��)Sź�sd36v� `p޹HC(y7:�D��G2��y�vږ��X2����kg������קj�*�,�U��g�՞�Q���т�������)�h��z��"��-!s�,H�����$JD6mã��?�-��o������}�	�4��Y�G�d��
�&R\*��������H��BP?��J�.˪@ؗ455�V@���~}�ũea]X�}�)8��Q��J(sf��y;2���0u8(�)��]���޻�4U�4���Eq�/�X9Y���2~=��E�GW�4�jm�F��s�}�^�m�8��II������h��|`��kF���W�K�> ��$��=C85��<Aa/�k����e��L�7�<<���9�抂�Iw �I2?޶M���p�w��^<3������h�":iyGE~��	*��)�F�$�@�pw+� z�=u�`?��sP�����=DQ34	x���M��lЄc�3��J#�oE9�� ��A^*�����aM�4G��Y��D�Z�ڶi:'j2�v�����feIgLx���N�= �z���)Ye���HN�1H�iQ;uGרS]N��Н.LXc;�K�� ^�3�̚�X�����`�3$�`�c� �T�E3��{$��	|��{w4-�k�	l��b_�b�� �L����r=�CW�ap�{����.�c8k}�?$c������KLY��ح��~�L+r�v�2v����e�kɢ�q7C�FV]d�d�vn��{N@����1z1m�~*��8�1�T�U���I��^B͗l�9�o�E������[j��O��Z�Ժ.��3��7(}�,5:i�i�����kUa�F�u���Ox��|��>ݖ�ҩ��E��Aͭ�~�-��&P�VǮj�n)��u趍n/<m���:�t_�I}�6��Z��B,{�D�{l����	(I��f�y���q�3DpIU�$@�����ǐ�΁	-��i��/K9?�Az��V�S��:Gi�wȼ*���ө[�٘R�����q$#��S��	�!�u$l��� _>s��������"��ͽ}Q�hǂj����4 ET�Ze_@T��0��=�~�τ�U(B=7��!He
��CZ`�/��ft��P�2{]�����XD�n���$OȐ�G�^h�Ly=&�zA[�5�Ӻb\M".2|����S3	P
5�QP�. �1:��p|Da0����0Zx�z#�}N;C��>��s��?��I��W�tY�5M���ɞj)ǿ�1�(�4�=Qҿ�WB����÷��I��~�5$L��c��|y@��ّu��r�V_"���S+"��d5��{�au����Y#g$�eWכ�8U�jN�V��<�����[,�X��e'`�ad��E�I9�'	�RFȲ�M����u�0��6�m��5������m��X�=��ķ7+{�q�=O|FI�"(k���Z`Xa�n�mk��}d��1��u�7	0+c-mi/\��J�!#jk> �^Bf�����]�C�^�h���1@�
�K�!���jO��mD��{x^�V�hK�z�#�L�(~Vp����`'�u\��f��E�@��ŧ�K��HG+#� �:��{������9�
��Y�7k%%��ƛmG׾�ꃧ8<�UM�Cж�������L�ҥ���Ӥ�0W�nq'~[�B��$9}˿��N�3�}i�#ih���O,��@E���>��H�H��|}_V1�/"�'P�1�νu�Qz��d�u�D����3���Ie���_D%�%C�t4}yJz�2"���EX1Ä��<����[kZn�OamD��<Bw�Xw'���d�tF@�/L�(�c7��E�g�BJ2l$v$�[.��(��
 �ס�#X�|�
����:�-�
�]J(���$֫j].
��/_���?y@�.�3�Z.���w|���W��x��X(�Ĭ's��?˩d�7�F���/kޏ���R!��������0���'-)P$Q�dCdT�䎯�t��,�&�.Uw������j(�0)�6�P+�'
�hO��?�-_�����.�?�N��b��s�kZ�B�%��뛪�����8Z0�#1�8k*-��Z;�@-�G��K��[��u�q�?M�����M�6,�]�&rm�����z�����H��X���zf\է��o��ωeK�!�[8�@"N��HU$�^���&�nY[�*�fDOe��k�Ǔ�C�vQ�J��KSL��ڹ���4����{���~V��Ca����,J�[�a�ye��K��6��s����P+��ä]c���m@���AA��j2<A���!l���:$p��Ǫ,�\9��"��J�,"Ng�z�j[A
�jƳ�S�pTÙ�t��Kh���?����7~�������#��7�9G�7R��w:×>���b�'��h�����m��Ϯ�:�o>\��(����A�o�H���
�=D鼉��]C�ڀe�Ym�����S��E�:9�,A�5��Y4��t�xXlB��b@^>%��-�ΦQ{]fJ�c���hVlF�(��0x	N�F��ү�#ɬ
깳e\8U��z<
Q�f2B����R 6���C������Чo�Ϝ��-ocX�0����{;10���%^�q\�w�6>=�+:�W��kGEgF[�����`:��e2���&e�����Ȥ I0_C��h�Z��Fꪼ�ߧ�����OGd6���d5���)�/U
\�Ӳ��[Gd�L�2�~���uS?pki#�a����ۏ����J1����E�v�����{�s!cu��I�||�a��$:��OW��'	ЍNn�q�^��z�=#-��/L����._u����p~���@C�b���T�	t�ҍ��0	��;��N���P�v�亇	�5�z1�[�&;S�jr���񿩛�G^7��XԜ����| 6�&�bƸ[��i�1�pe:[]8���}�y��a0Ă^������b�HV$l3�91�����I�6��� �,ϥ�
����U�k2+`�����"$�I��+�&Ŕ���J�1;�{d�[!Nh0�&h
���;�#�Úi���b�Qr>��0C5��ܠ �H����R�V�8�x|[���<*���%��R�$�`XE��TD�rTYu(�ۖղ��#�4C_�,舢� �j@EJ��˯ψ�Ϡ 0�dg$,���{�h��X[k�@�	e��'�k��X+4S����P�P\?6UKՑ���#�.,
XC����dZvB�ꮩ�5��0CPLު�ކ�'��袱Ov��P�a��+�؈��KXU���ۭ`	�sI@��Ԅ*b��fl���?u��ǣd��s�Ƿ�˅��4��{�8��.�5	���q \�����M�����,�q�k���8C���#��ؾ^���U��֎�P�6���"=�r�S=
�jI��'cO+��UF���:	���P!L���� 2�1�9�� ��P�A̠�Ɇ!�g:1ڟ�T�Iɺ����H��󆎈��N��4�2Y`4+t��S]ç���j���E���p1���!��pCaў.ّ��xf��m|%R��䍖��6�:G��P��F	�h�=�DP�}���q�.�ۯ��v���� �������'m��꜐����ǚzP�#Յ��N�/wS�ߎ_���i�4٬A��Ay���JwEۘ��S��Y���o��̰L��_\,}X3nG*�'��(rv6�TҢ_�K�.����׍���Y�;wX{��eQ?&��"ؖ�����I��Hgl���=�=�r��2����D����N�~Ә�G�����@�A�1�<��9q�u����,�i�CI�qab�����v�P�<�����F��O �B'|�C���R��-y��%a��&>$���>���3D���⦁���닌܅3�О�r0�Zn| L	�˩��k�@��u�8�5!�8�v�Q��*6o�ђ�����mZ���<�^����Q�I��+ȹ{����8�H��T�_�<�i	T���e^L�!̲E�WS���ۘ=� �Lb:�]/X�Yb�U����5��}m�C�^�}��F���{y��}J�!�wI��rk�{��#�!1�^r��^7;*8�O��D�'���d�#{Cp��)zeZcC?P���5�m�z�w��,��Œb82ݘ�Hc�&3jܐ�l�~��A�\5t>�Ѽ:_�g#��V���p�Ŷw�����5+�U�`D�^ۏ'mꇵE�)��Z��G8g �0��7A�|��v�o��aYh�j]����o�����f��������X��:�wI���%A��6 �$ؗ��S�U�ؾ�S?��8���lv0�e�k{?H6�-&��r��A�z�kB���@�$@ %��ّ�n����0�u�D�� �zCi�0B�Q��d,;lc����X�`�^J�Y-nZ�z��Eo)������W�Y��aF����9cR�%���p"(0̼�����m�.�dʚ���	����p�^��
-)?i���\��iErrqTxV���Ol�U�c��º����f���XS���XS���Y55B��do�2�[|�l�P�C�&u��b+P�doYϡ���B��b������Qu�r ����	��=�2���;)��q}�?�ϝ�gX�O���I��ݚ��Dx�6O�[RG'���Wu���f�� ����W�~ɡ�cq~ �U{jU���ڬ{�C_�H����R,}wM���fkR�-���7��`_��s�,j���[m�"�U�K<<�������S��*8�QcC^!�-k��	+@���*����*e��;D4"r��.�Wg>��!߆x������%��S�h�c�i�� �sw2ƺ���Q���,T��o������Pb��i+��j��~��� T�O�ٺC�G�v�D��KՌ#a�1Iޮ�s�I>��V'�4��	ԕ:�Ɇ����U�uq�e�5"���O����o^���yZ�#u������s�Vdz��W�@V4q0ҏ$e���&���]縬˻|�1蔲T���΋��#�qM�\�A^��'�#���F�#IN�E��/�	yѻ����p�$OBa����f�3/DK7R_ 4K+��*ũ��jEV���e���b%H
���%;��tB�'��[�ޮU�s�U��"��'��G�8JſB���l��U�^*��]� 3.���Z9��������U�B5���Xʯ
�z��2�P�R�Ys�Xr�g�V�C��5,K��G"*[�@#���L�"
36E7۾kB<{��`%�k4n�b򓡸���-������o" ���v-�g"_��"m��]�t�:N���b^���(}�����O'E.�z�^�k_��:�������̀�ɲ��'��$�M�[�}8g��O��,i�(=�]J=��w��&���̅�Γ����@@b�8��2����e	�^vAX�#"<�������U'�r�WR:Ng�	G�4�"-��#y��#��r�V�"�)4R����7�{&&���R�<�8�tv�!��?���mh';*��X��=[hp�B�x�q	{ς�E�K���fř�.j�R�F�cX@`Q��>���;&�̶�xa�!#��%�YН3޼̠Շ>@�)Y!j��%�T��8��:�I�s�S*(.�,�?����/X���e�Ds|��ʳϽg��:��pt�c����ZE�l|�qi�"��eQ�g�١|>��MNm�,�^-=[B�P?4Ϗ����M�-��w�ŵ��.�h�0k�����zR6�h�7�A�OD��w���f��l������/�Q<��Fd��l����V�2�	������̓�����,5���������_�m9q�h�^*��y`ue&�����`���@V8�B[�	Z=�cQZC�~�����g��ʼq�	
�����3٧|�����7I�%�,Y2Ηu�)�.�:b�$�h�_�N��z=#�O�L�P.��>��|���^kk�4���H�r2r�������S9K�s�.� ��]�N�#
�$:.�\���*]79喒�i�0��(�_�VgG˧�n%\�r�^�'+�1������~�y|1��y�*���ܼ@�A�����Ȍ�Ul?x6��}�{����^UXe�~����F����<�����'�n�6�{R��|S�*�<�;��	�Xz@M��v��+��(Hcw��4}B.�9�g�(�O*�,����aW�����I.ۖH0��h�U~t���XlxVHYEB    964e    1150ҭ&9g/����l7�t��.^�z�~s���Y�8|���:�m�&�C�Z�bՍ�Y�w&Ph	��n���=t&~O B{O��`�֌%�v���)b��6��Tr7Ǯ\vK�F��qO'���|��CP3y����؜��)W�������)c�V�@PM�ߧ��Mhݧi��@^���\p�TP�t�s;ȴ�����P㇁'�8|&Vҟ&SU�j���h5�\����j��mR�;�[5���E�
d�4�m v���B���JXt*r-�������<����<tXG�*�m�R�yJ���n���`��A�D�����m/}��8�����j}��[�|
�J��x��w��D>�#�8�Y;4;Xa���y`]����q5W8��SBd~̵N:�"ڇ����Js���&X��Z9��%|U�pP�!��!��mz�߫bsY���r�[

+�nE-�?Ş%����'Q����a���--:����~1{�!x}�h�Β(M��ǈ�T���~��X�*�J�7FR�p=��ܜ��/�.q�e�	����o�s�b�H7�׻/d�W�%6�a��"E�Eٞ��a�t��Z�iT'B`}യ*g�MH�ӷ�.r-o%�lw�"�D��5���W��V���Sɗ�.���2��TAE���%�����b; ң`�ŲB�������y!OO�6l��\%�fOg�Z)�+��n{A@�G5>e�T���xwh��!~��?���h!佰Q���`9W#�\.��{�d@�Z#m�8�E>K�+cy+�-�"��O�t��|)��I0����9*ն���HVK;�/��
��Q;{o�'eI�Q����b�� �ݯ0.����������������H?��?�����c;+�M��*̸�|U����(ȓX ����O�����*��;3�q�}�	��kʠ�������r{�DbD�ʍ�f�3� H�� jnb2O�@��mK���ޑ�]\~��H�X[2J��.�<|�O I<�FQ�e�;�~^���a��<6�|��bF�V������m���� � z4��R������4�P8~�+��ej�C֔GI.|����E�<g��+�|-�_���s���X�G�2�?�>+�f��(�O�tGɳDK�9Z�R~���JC)���M��C�����4d-CEswnqZb�_����/͏g�ʋ�{r�z�kBw.��u�����s����ht(V��~Ad����g�����p���
�̱8Ӈ3.�Ѝ%'@�a>N�Fa�U�v'�E�	PSN+U�xU��Ҷ�;;B'`�����c
��\.�{�{P�	V��H�^�;V�#�MZ�R��K����ose#t��ib8>�nOLF�84/놼<.��d� �Ň_I}��
����^łX=Q�  K��D�tٷk}���}�38Hag�u=	� ���?�0f�٬Ւ�Օr�
GT��Ǿ�5�ZfN�5�sKY���'�͘�n�ŭʕ����	b�������J���ԅנ�8k�{������ݎnTI��l�Uy��oɄ!\/g:�3�+6C��� ��F�c���l�?3�Y٭ͫ������a �VkvG�QY��_�����3]"s�YG�7҈������Z�=�ΊQY v�%��ms������{Z3f��8]%3��_������[d7���f�E��$����Ջ�9�\����k4p��Bm�8��W�űG.A5G���4R�eme�0\�0+�|��F딹�}."��Cg�jQlF��r6	bh��X}�qǵw�S2*��o:<� ����Qg��|�bY�{�u.���<���Z���~��8	�$�xk�1^Й!k/���:.�?���sx�$8@���]1�����NEܖnݍa�
��Z��z�æ����t��2�z�Z87�N��r	r����wM`����"�pM*�\�z�n���U�I��w�%�A!��W�}�9�n1^�۶j�UE8����� Yq�%�$m�o�5���� ƾ�IC����������A�,<7�?ܰ>�W]ś���6̖ m��H��ۥ�1j��.��Tg���{eTw�F=������w�oWo��ן1��쾌�N�c�3Gx��v����f�B���	�fqg%2���O(�Q�N���sT� �,��~[�
+F>=',g4��	���?�=ؖ|����"��m������kl�n:1_��@�ߢ>39i��m,�Nt4��4A��"N)��XZ�̍�`Dω���D���AX��<>j ��A&�5�&��+l��3�u'�~R�l@��W�FWsL|=��$<JeQ
Y�5Eq�q�^*U�x�B1�B�&IBK�N�\������g���=)����6+e^dz�Z��B�w$D́֧[�y�	��z�e����g�A�Z��� J�<���k(1��:R�㌓M��ߓ��>&u\:eL���"�Wq{�:����l\1L���9ӣ�=>�����J�m7�����(G6A�B�& ��&x��JQ��輟�����z�Q+@8��<�b$�S�h���Sh�j�~�m�/G~�*�M�-�h0~|��Iܶ;��\��>��W�f�"p�.�[.ln�ey�s ���^�`��ǘ�[(�uSX[�"it�x���,r� ���Y˰|�Q茟�N{W<�7(�֐%
%K֫^��VM+���_.�e˺8/��k#SA|ÄE~�#{E�)�����Zߚ�r�N.)nmS�����!�����-�bJ������g.��-]�X9i�����bc�DB�q	ļw*�a��zN���y�e�+�L3���S��u�����*�3��eA	w�+;6�aY��6�=t�Z��-��7���9�:�U)U�[�R����L%�����Ǖq0y��O�⢽8��׻7��pV��v1��y��;�!� �G>���b�~��]#U�I��˃a�*�'�K�"�GM7T;z���E5<�%�o$!�a�O03���S5A���'�&bT0i2>#���S_]�˓GBO#���H��K�U��?x�� �)�T�7N�L����hu��(~ ֕������I�� ��f�G��n�-$��!I�0��Q��;!YYLԁ����Z������4�!I�9iy��`g��qR��i�v�5��y� Ȍ+�����𶟪��w���䍥�~
m���%��2ɘ�WR=�VM_�1Қ�Ҩ��BMWp#���VvK�>&�ALd0�L���/2�6�'��G�ix"p�D4�p�J������Φ��YR%0/p[�)6�>~b�\lE!�?��&������cu1E]Tq0�MQ���^�n8�a�D�Y�����Rϭ��h��Ӈ#
��9="��;�Q���������/�?��v�+۔�%�Ru����F8�V��02i(�q��h���<z�s�Y�d6���r���6Qt�%���ٷ�%����ф�������SH4�4�ԎEI�S%x0v�~:�<s�h��o�J�8Z`;(�Pkk�gx�)A�}],��g�	I��g�u_�����N��此���neD���/fl\DxƠ}CR"��H�L���v�n���&��r|�a�(�⥽��=&(V�t������^����Ǻv�?��7��W�a�7JD��e||j�=ُ�G�m�l7K�d���-h˫�pyu8*u��HM���:�J] 7�@`:n@�U��O��Ma�����<"f�
@Ħ'�S��)H}9����0. �ը�̸��$o���jD'<�m�o�W�]R0  w�[�5�J�.�&���37�x
��M���ܵ}�p8 �\����x=�l$���@m��[�g�o��x�<_��V�����K���宖��7l"����t0 yq�����¢7��#RKH�ms�;zr?�k��6�}�ّ����!��D�:v�&g����Т8~����D��g�~�����5מM�3I���,��kpǠ=�L�Y�&�lk�1�Mt�+�ַft�u9�ռA�`E��O��j�W�L�})P��)�p�ǀ���R�����I���T+�����ʽ�( �?*�2��i�f��_50����hHj�'�6�q .������x������A�=^�ХY��
��H��b���Z{�E7n��P6��24�5�}�{} l�<[��R��8��������X���� g �Ux�9��Kƴ�q�ǵ���/�b>���8�m�#D�B�3r%��O0����W�h
.冭O���M��O��3�Jvs��e�'�l����e�Y��bF��5�qm��v��!��bk�V*͍E���2�~$�����\��Ay@f�<