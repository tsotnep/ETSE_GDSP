XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���O���>� O̡ZT�m��|Wl��X%dԔ�>�Of��O��G̷㗓��	J�'[v@ڧ~V2�Q0�Z "��o�K$fu�|jk���p�촜�6��in�,ܮ�_٪�#('2P�A�[j����HNj#�у��'Vh�ik�N����n�g鷺�0jO	Lp�U���E���a�B�ߛ��j���T۔7���ص��A�B���pb��c���0�pc��ٵ�ް�r�[=���3F�e�﯎����Ŧm�����]�B�[
M`�Be_N݂�hK�x���I�H)�m=@X�m�y�pI5D��E����D��I�v|�0�ܬ(���+��Ƃ�s�k�_��o %���9=O�����B�C�b����$�j�&9�8�讈m51�b��W��"t����`��t�W��ְg�o�Zl�N�t�9b���5�����pϺ4�y��Xy��� ��w��*£FB}5�P1�C�~e�'��V7Ú�څ��N���6�|pNd��-S颌<R�����.�l�Ĉ�P5��J*�2�ѝh��\�m\�S�G�7�9��N/��=���wY�}�b����ǋE�|G��Q+'�:��G�-�A��sġw{���ڂO~���̄SOY�]��.����_���۵@n�Q�
��dJgW�#�<�y`�u��G:n+��h��t�7Y��VX#M�<��}G�Y�!�o@1?p��?���7�gOwԂ�kv���cn�&)�@�x�s"�z�>��XlxVHYEB    fa00    29501_c׵�>��������"j����(���$��n=#��>�}��.ɣ��(*���ru�x��}�:p'�Ri�����b��i%����2ƙg=�z.1),E����jۋ9!#{�:��p(P�$=�L-ţ�J*�4�v�a)�)3�]xW�.��(4�j�WQE�V��M�3�&�jj����u���U�7���o�� ��J�����֪��K��!�:g+�3���l��N9��j'�d� ���~�H���d�m5̢�4��h��^7�x�qV6U)
�տmގ��G�h.�(<�:�GH˜d,���&E������<�d��.����ØT����geR:,� h���N�p�$1k�B_L���.��|��	�*�j#HP��I�acTD^����=� E��h�� R�������W��)+��=c��?���4%W�h~/�Z���[��^��#��o�56}��|��­Đt�[HRR�
�) �#�-T�� �@HL�v���%�4	����L�/f���P,=��0�g�C�0���)����>�����ռ�9��%
�fe�-��z����	ˊq�UL�^�r� ��	���㏁!���XI��21�*Jr�lL7��F��2��}a�M������
j\�^�1���̋���}1�JH��M���Or>skNx����[�o�v�h	b�Y���(4[A�������/]��?[k]�Q�H�`:�G�3I��m0��&���(�AR���5�uv��L�v|���
��j^��q�<)���J+�^�+S��-��8����nD��8��t�� �R?�aZ��2��fR����jf�1�tDBՆ��zM-N+�
�'Fcm4u�(�b@���	~n5��}���l;J�<=X�AO�m~�*�u�net�u �i�)8��h!�J=�QнY�c��O��nҬ�y 3������"0�,����Ơ�X֏�Y�������)@!���c�߾A�V���Wl���ii���U��9B����0"��	���A{8ͷ�,��(iʖ.�v�K�g���zX���"�uڍ�B�6�j��������mQ���g�wBs�!�('���1�fH�Wsp��E7��	!�.�5,W�e[�ո�?���������W��j�/�X@=��Z �5�q=�������w5FK}�!�ÂE�_�W��OSpe&�Ί!�y44�wq�A���+�T�r3�g���׊�@s/E�^w����@H�����g��R�z��\6��oU(-����D�rd��&�Vfdp��� v�N,��Ȁ��$_n���� ���3%?���?���#�D���r(Z�[�`�V�*�� �?��O#�Y����g+0��Y�U+-��@�눼b�u4��`n�8uϨ,�Tp��U�8�_�;�9�H����|����Z/��Θn�,f N�1����\r$�2��`���1޲hw<87���B�s.�[�(����#����9妯�S�������m����q�8p�Oo��MY�md���]_�=}�;Q���.ũ�5#\;�S_��y�{��WΥ_�i'yv���z&�W=x<�����O�	E�/fx�n�t&��mn���#9�Q)_��3��t���Ж���AO��R`n��wC��������� _Xx
�����3(���&A:�ʮ�Il��X��/���h�^��TO��E�܁	@e@r�	�.����G��ٛyM&�-�2�����XJ翕�����nc�������(��D3�OS����z�v�x�讎����9o�T�s�#A��ꧪ���1��';@�J�^V-�/Hi�`�Ռ��c��R^`����j܁�֮w@�b���� � Lq�U�d�y��F̯.S�_�LeCg�d֮�O�_���{���Asm�4�/\\ � �G�8����������W:�r��P��חCV��9�~��S'���lA�/4�_��ɃT�9��G��u�t6��LΗ�������	��.� o.����V,f>l��Uz^�Ҧ3�^���E�����ɿ������~��7w4w��W��n��X�_Q�푎���(�O�����Nbf��1�gv�	|am�\|&*~c6�m]ٰF�Gg��Lȼ{H���ܮ��Ƒv�?�a�li6C��uڀ	�г�B�MW���$�6��A�R��r)>@�+��m���'ӌbq<z������\�W)��� �^r������E��4�#T�u����8�K�1����J(�AdJ2�=\[������Q�Rg|��M[�X*a���B�B�V�Q�}�Vp���*e��טJ	��v/+��f�>��Ǝ{;�&� �-MzQ�����9^���a�Gz;̣e�,���������؇��?�\[*�ʉJ�����V0�*�|�w�J�(�f+�(Ta	�T �|�j�����T���ʰ�£�,>9�5�#�>��8&�k+?���t���Ʊ�d�+(���ÊԼ# {"���i�����g$�=�- ڔ"��1�a[oJ�݂�c�)1v�d��2���ݛ4[���~��n�{���+�'0�#�����EQ5�Y��4�Fg󀅝� *~��7��		�OL�(�<r09~���+��{���Z+R��}w���g�Qo˫]��;ek��
��?�T�ߺ�'
�w��R3����TH�Y]��ros��V��v���s�:��R�~O�hKH��{�7$e����nE��D����fc�PI�А�����P��0:D��(�^�l�E�sk{�$V��W@�~~���d�� �����4io����zHd�[($�\�2A�ȸq�c���@����n�gi��dvc���Xl�|�i����{�����	����|�����e�O?a��P_����ʧ2b��z�%G�)�5�2���Dx�ź��mM�oUۮ��	nw����k��ٴ��uM���-��U_i'�O�ػ'�'Cx���\?��E0I�oQ�w��jH����U�o ;_q�-XkT[�p��L��?w���/�88�/�i�pؓ���u��u�������<��D-T���Wb� ��Vᡞ�c�o��K����-�E]���QRs3>��?ϡCfܕ!nC>�����f8�W���xc���Dli'"��enz��=W��'�/��NʫtU׳����fN�`~�M۵4N ���%b���SyK���:�I���c^�.>�%~M4O���=�љ�ޓ0�9�ZMD��
�4GC��J�c�΄>%���*�zͮȁZ�t�|�)��+��u���8&3��9%��|��wF���}.I:���2%Rz���$q���?bz�޳�g��1�'hx|��sV�NX��'5�G�mȔ��x逺�
��	ͮlc0Y�VM��e����}Qz���5��ݨQq���TU�Ո��z��6z�T����ͷ2��O��M�
�����b!����M��V�����0��9�c�������A��r�� �dn+�&m�[=���C�	\!�q�3ȗ�5 ���I}��\'��iɺ��9�c���Q$��JJ"o��Q�YZ�;��|L���]�_x���ӷݺ�R:�����@���J�?��/��Y�~$i�æ��'�lj�-U kˡ�{�Z�?+	n7N(n��<�U���q~�r#\�`�lmb��ZMo(J��������@躬���L|7�Gp��#��xIWuz�%g.�f͙�e�aFr�,��r�]�Y@ڋ5heq�(��h��7��$q審y�d���MC��f��9t�=Xcvh�`�%�:�Hvі �����%��H�X�7�:�IS;�Az3�>��������.�	�����|<+I�IV�����OR�`��!�,�$"qK��"�n㕚�J�
��Q�_�S�L�E^�1�ճ���� }�Ap�Qk���8�
�t�^�9�D"��:]��˚~����sB����Y]��`
�ѵ��h!�M�l:Oֆ�Qa5�`/�h�{kP��*�:d����U�>՚sᣖ�x��t4��y�	���h��� ���&bo0d��<)=\N鳑L��Y�\��y(׈��}���ىV�Ƿy��5#����5g�?k�y1zc ����P�6d����i˜E3��˭��7ej�wF�T�8�4O�rmt�ݭ��W�mp&<��z�p$WV�=D��w�����Y6ux�s���T��OJ#�w+J��`vm$T�e�8E�>�HD�pz�3E�W	k��:�W�X�����[m{?�����b�@d)�C��̏�,��
t��О��	�KH$��Hd��T�e���	Σ]��|�޴�4#���x%#{Σ�i�!ԪFĤ�QA%��pmY�"#�ҟ�_��2�.X��9��f+�0���K�S#�	�M`ߒ�[�X���jf��)H ��ۿ4�W A:�vI���_�g����r�˽l��������b� .�Ղ��T�5ζ�؋��z$�j�P���B3C���*��'wia�iip|
?�p��jh���Q� �k'c�o�� �CG��O-r��z��H��!a]�^���m�����F[5�
�1K��mRX1�KI~�n�'M�@nAS��bs3�ƒۣoom�R���DAA ��|��HN�ƽ�'"[��P�Ui����0������)����ݹ�-,M

����[-IM�m�c%�@�Hb��3N�g�x_��S�9̹�v׍8��vY��kx�\ ����*k�,��a�x�K��tA�fB�i���ͣ��%�~F].^^A��3�jga�n��E.O���8���ܡX��i8�ux�O�aW�{_�1fOS����n7"���GN�_/h�I���"��xͥ� �n(�\��]�<�
V��^$&q(NNoO�C�Wv�[W(�E1��X��v_/��ʉ�u^���͚7~�ڙ=O
�Bu���}��~��/Gt�$���]�����\n�3�M�z`yʿ-,㐕�dwz]��X���f��w���:B����i�1Xi���L��D97%����L�h��w��?xP�G�p��'+��xP��9ѹ�&T��;����a��V���� yN��+g�]~NA[G�ɑ��3�śRWN���sؓ�e�E��N�ӿ`p,Z����7弇\s?�Ꞹ �t�ug�o���-����	�3�<8(l���������̜ޱ>�O�+Bp:ǆ��"ȒriS���o�BcL�&���HΈH��\�E�������"ت`�R�c�fer� �\5��
�T6���m}έ�y	���z`M�0�e8���گ�aǢ6 ^��{8G�:���׏P�p/N�$�NH�{p����u��S��GɬBrY�\T�o�KHS�td�vX�@����f�WxM���F�%�v� Hd� R���76g�9��(�&]��˫��sv7D=&ޘM>��W��P���]V}�NZwC�v�SZ�=����'S��)	x�_lP�ﻃ���ho�t#�6 ��i��܂��.r]%F�%P��zϧ�!#��TO�H	�����Ӳ�y���b~���;�Ɠ�h�bLأI����8�{9zujp�Ϡg�����G��x>Gbv��ד�L\\���0W�|m{�Ìf�H�[�K��?�]�/�$@B�Ru���B�4����ϒ�)4pg�-�N�ҫ���Mf��km�n;c`:5�#%���G�T�5 ��fKS�~�^=�e8[�f��u\'^�/�{>D�03Z!�!���l���rH��.J3V2��� 7�ī/w W0Km�*�M�!,b��)Ë{��sd]�ܗ�,֏���>3P
�09��T8^IC�S�(Ŋ��D�#�	��@��v��� �wӊa��֟��A
���@�}���:�����)pn������ai.T�����0�v:0*�NN&�7!@C�:��s�d�ѷ�C�5���عA�AƵ�nԫ3g�(
��ա�i_x:ip����H��)�(��f�ڕ�у�>�'&7���HE(y�iyg�h9y۟�)2�C��v_��:�~z��H�5��"s,k�S:0YY���d���Q*z`�fbR�!J��W9�xC�|ʫ&-]�j7p��㢙�f]I����� rPed�v��U�6l~
)u�}mm��Y��S��dS���S�,��!��˭�ߢ�p��b���yſ_��k��|=�[�L�7�?�9#l���P�z5g�h @�����]Тa�u��~�a�y]�����d>�&:�R#�2���چ�<��0�$b�#s3�QlW���s!����g�Hz}���7�C�	a�u'E�L�Z]o�mT��N��K�|�M���2��@8���)�5!BBZ=�sݞ駉�Lf(��؋�G���f4�Ԟmegy���+�y�����o���r*~��t�20ҩ���yNg�qS�L$����H
<�HD�ˤ\�DJ�E�-�`�XTi�*��kk�Su#�E��nZ]I�Ps�;K�-��r�m)��f_�ށ	p2Tp�YD�-ݦ�1R)q(�k+gs�B́ z�6`ŋF��2w�`se������d_Z�����0�w�uC������IU�ph�W����u��B
�g7SFQ$xi�����4��O�?��ngs^�~#N�^�z�{|�RȒ ��)"d�w����+�z��Pr���{!s��)��I�B�Z�'c�D��Wp�M���$�cL(2x�_kFNg]�@\�z����ߔ�D VL5�\}�<�<Y�p�4��ie<)з�S~����!Sz�\������lV���eα �*%dI�hg�?M����X�����j�n�I���7Ir�t���(�U�s��ڀK1ȡ�J�����z�����cW��Ű<TM7,c�5r\T���>�����W�רK̈�չ1O�[�T�ru�p0s��8+�CN��;ƈ@�VI����/��=�H��q�&9
�/�ŪQ����x~�%���,1��	-{��&��0U��w�f�{B���	C�V��D����_�w��]��'R�w1a/���xP���5�B=Q!�!�?;�����4a���"9�z�X��,����m~H��LX��)�Ȱ#8	��>:~H94>������K����Z���F��\�3`=�'���7w8�F� ��+�(�4��G�l���m�r��Q~����3�pq�w7�jƊ�Uv�4?n���g�cQ\�[?	��Q!@+��y�V��c��,���`a��oF�Ch�7����R�����Ew�N`��h��֒ϧF1��^ΐ>���v�Ci3�;Խ"H���}�O �"�[L�'����VEq4����� ��s���?�ך���K6�Y��л�� ��ߚ�Z���%-��S)����mj'�d�4� ^+z�@G��G�#V��ǣ�[�-zQ�q&T�5��2�|Q�'G�G�L�����"����-�a���W�t3B��?,*�W���S���M {V$���3�ܒH)��#$�%'�����/�0S�?��{����k�=t0.O%���#�8��q�1�b��R�t=\gY�6�
l8N��bsǹ���)�k���h�޲��贤0W�{ɦ�@\��͑4v�,�v���p�����cwm�Z��(����+�����ڳ�����h��m�E*���z5!Q��CN�,�jg��O�\���Ǡ��e�ut����M�Yہ��b�����a��<�.��ԅ�`p��{���w�T�}w�+�tS;ȥZT�Pmt���k�ؠ�rK(A�B'�����3���=+d~GK���O2����;�d̔'��꺀%a��
��<�v��>�:B�и;ףh�ٱT������L�c�ǈdA�18XJ=y����:Zԝ3���m+R��Z~kD�冄x�h��G�%��Tt�qN�h�׭��[�)��OA��[��i�f�K�.��b����&Bίd�Vkj�'��\��*�_���ܺ`I��t��W�Ln��9���s�'���wT�rw̭����I9r��QW��w�����#��~N�}d����j&;L�@k��"����/h.��"�����࿇A�.�4���;|��h���$�d�䦿��D6Z~Ah�Oh��ω���c���x�*GY	'�B�9�=?�ʖ�RF�s3|`�<�J��W	R?3m@�vw,��~J���wv��-c��cQa0�H���=�i��q��͜c&]��d0�{�[)*2z��(��5���as?y�v��uL���U�-<D��:= oO��0/����/p�iI�د���b#빞����$����ׯ~&������Yx�m�u��/J��#Bp�F�ۑz���K��$*|UR#�S�FuvI��U+Q&o��%qIn��ߪt��ܦ2�E~��e�"��;��*�L{a�ܙRIv�(aH1�.i��X��Fs�۟�zE±D���?�@%���~��e��b��H|~���~k��JD��7|�UdV�5�X�����I׈�dѴ�Lմ@870F�cv��.ef���Y��Ơ
�q/���H{Q�F�mq2�c�!@q������2��2grF�\�6O2($��_M���*���v�Y�H���A*���PI�=ϗ{����Q�g�أ���y]�����b�X�M��0���Ӹ�Or�ܳs�DCZ�N��tyc�i��/V�.�w^Wg��[�&�V]n�2V��љ�O�d���7�B���8oR]R��q��K�lR�^h��!��"
/�0׵�o}t�u���ۛOf��d�l�[�y[[����zv�./^r�3��p��w��=�*�w�:ё�v�39��h�����1AU��j1ǁ4����<K0M�j֘ {v�U�g�����f%񍉵����1�f��ш|�;��*���Rx]�ۡ��u$Qx��u�d�
��P}��~?���W/i ��(�����X���7��ʝ��"��WUg&՞yQ�7`��wt����%��Щ��ձ.��^7{@?�$}g(�?�Cr�!�Ae���A�ܕ�T�W�q��N.Op�Q���B0Ĳ��D�.�$@��1�8��ܻM�o�-�E��l�Ec85Y��@�V����OQPxI|4I�+Z��j�(k�i��m��7=3�V�΀/�o���cs��yo游:P�7!�H��;�y�v m�z&bz�Iő�tLO��Z���\H!io���iS,��b���R����ʕ�$3�z4������8�Wںbm�Z�*ו��q�lc��'���8�fǓ�S��� g)��s���ac��k�_8��G��Ԯ�9�����Q�x|n]�B�
z���>�`Fɲ���g7ԗ��7�Qpیwq����Ξ��<�'�.����牧1���3l���s�1�_��T�!g�DZ�\Y�Ia ����d=�VZ%KOՖ�!\	�˶�|�q����A;��Ed%�"���[8�(-F��
��k^A��;�o�P��MGܴ���?�l�܃Q��v�_"���/=�V2q`��-̤�,:��l, M��T�~S9ٙ��fǆ�}r�=��|ή��5٠q��р���Foہ��f�.�µ��گ�C��"�>Yh���ˏ�u�Q�ʉQN��1��q¾���eC�z��ߧ�2"Q�V��ɍ�g�!���.��U�
�K�`�^\��2�[Àu�A�`�^�É9L*7W�3��h�ܾ=��/Ξ	6P��/pΜb&A���4����l��O�vfKÚ�_Շ%����?�Go����2��W�Q���#��2"8���OC���s��0FbK/s*l����ǻ/�6� �0�����'1<��J�~�ؔ���������	�(]0�HyӚ{�߳���I�DrB�����Y�t�2xb��r�+u�
x_�ւ��/Vb�Օ�R��`�t����Ɍ�iCنW�}v}qLN���P�SF5O'�[ieE��~�B��S�ď{4� .�sM	N�,�p�/$Z���]�2��e�)��7���"��d曐�{�?Xi��c^A����Y���e�k�x߈)��G/���E����_��C�=����|x������ϔ9��TzNQ�㾤���4�S��8�0ͫ:ܲ���c
����Vx�<����S�G:@f�y�|�m���"���u��K%�[*�~W��^=Oy	v�n�ȵ����"ʪ<��Ҭ�/Zqw���a�������=o�Em��H�1��wP��"��OwP�����G�+{Zl�w��.���'����6�Q��)��J����?}v2��o��QRx�AE�j�?�XlxVHYEB    fa00    1e30�aR��y}H,��]�AZ�ʒ�O�K�J�3�g�>��'11{f�Y�8�X��و4u2���5ϣ_���,�8���6�� d.�ᖥ��6��jU�9{<ܧ����~�h8�_dJ�ϥ����'FD���F�/�w~�H�^G�=4�bҔc�W"V�o��L'D�KlM�rÍq��3���xo� 6x��UGh�����4㵩+z!:F���	I�������m�P�B���� T�XɊ�����>�DY�ν`^h��?{��tP�
Q��cah���\�"�'
`n�R59�� �VORj��9���_�W5��d��O�G�J��j-��g@��.㛬�
<.���M[��y"� �J��
���ք��mrp����+i�ل��d��U�W��|�,��H?��i�����!��k�M�l���%|��|V(�9�ܻ�y��sh���l̰�pbw��G�%>+�X:�e�n�&K����	}�B6�% ��6��[�;].�f���ƣ�et�oa�܇��*?���',�����<��L�E/Tvg+Æ
�����:"�(�lv����}�C4#�� ��� br&�#v*c�	��]�/������xhL�8ᒱ��T+ �Y��R]�q�DQC�)p�
y˲;a+f��~�dmr�=�MJX��ۂ��B�Q�"*%�n"T�1����@�*S��Ԡ(w�.��^bD#�����7��f�_�$�Lȕ+z1��j�Q��N ��.�z|m�Y�BYPyc~O��+b6��
��\��w��4F[���r�H�rg���47�K�wڈ��1�.W��r3�KPF�ԡ�z���
9�|z�H?Xa�/�g�_ES/��=իx�O�]���U�g���{\���@Î�����m��2!�ˍEs�Up������s=��P2i���Ϳ�{�:c_m%�!�5gU{�O3�RK[qg>�a��^�J��&�HPކuI�^PU�?8*��x��R������s!uH��Hl-�
Y� �m����g��5=�>@���+�d�)ZH����HbY������*cY!��zwX�?�Yq[��g=K��7���w����0�%oL�y95�(K�-u��/�Ζ����j�X���P���&b0�	2�_�+�?�f���=��	B��������׬]�jP�����{W;߶���¼�6�I)�iA6�'6@��	�"�f�濩+�B-u8+%����_闖�K+b�4r�I�vɒ~��݈	�h_y�`	%\�~�_v�`O����?1c�������$��X��Ī��Ŭ�0})S<T)T���C0%A�0Y��(�[*.	�U���4jLg�-4��Ö4ǂԳ#`�:Fa�b�!aL�?��&x��	�ƺ(�Ia*�����S.A�nVW�<9|=R}!Q��������~E��g��h=7܃~_��s-�s.��Sa^��6�������ݰJRS�l�L��0x��o��<�T�E S�]wu&+������O�@h�j�F�N�]�q����=��>��fW6�s��-a>����E���4�Yy5�t��zH
T��ư�r3edug�@-��E?��p� 	�?��k�\-:���qq�W���L�֎o���*���VPh}7hZ0�O�u.�����c�%�iF�.�tVAE��c<<3��A��=o�n�59�B�����O���B�m4o���UFJ�j���k��{��J��m���>��� O�q�IQ6l�W����H�e�Isg-Z�d��p�Ǭ��SC����+�G�V��ƴ�N��Fz�B}��̳��-�R{�O�Qj�,R�p��M1�2f7�G���L��?,1���s�ne� ����Ӑ)���*�v�1��[���v~���!�R%}\��G���,*�C��K��XO|�^�y7�E9ͤ�F�����M̒ĥ4�/,�PZRm�M2@���������nf�HbES��@%	b��j��e�4��F�F�G
(r3����v���%�[bN�8-:v�`��K*�H�3�\��\K_2� ��c��zڋ߽e��Szh�-.b��2M��Z����4�7�\�KÛ��"l���%I)�I���IZP���e��w"1���){�~���"�@���﷉ĵ�Dvi7x*�ˁz9NO��,���[���r�:!�:�"3и̽}4Tر[�&?�^5	�>��:U�s1�dG����������S�6{��K'���21�W-><냼e��UIQ7W�6V�7�qv�>DS�U��)�#��[|3O&��Pl�Ml�����"0�=����8h?s�w�����<7�mN�G�����s��i"��짌-)r���Jr1��%/���^߻�up��	8b��[���c����Vެ��Y�m�'�&�`O�ӵ��������p=8҇�NwL���o���*6w�}_��{{�k�P�R�9�f���6�,��z���:u�)ȋ\�	�
�:ǉ����ְTV��9�/�'�Ҭ���b��R��'7l�
g��`�s�ǩڠ\v�e�����<��eD�_)~ܬ�T�a�"ďD��[��;_�mH��mgN�oy��/���-!�0��-���>��3)e���s�R70r�ӆ����?Wv����o��D���4Х +1P�,s�`x:�&���O}��'�}��mW lK�䬚�B�ٔr���A���℠�#2�0c		'ک��Ț�iEz�"�~��{�D�6Y$�1�� ��cɃ�uU���$�/��D�w�0GU��S�������AI��[�p��N�ˢ~M$�[L�6�'���%������TWL���[z�Јa�R6��B$>����kmz�4�JF&X�EZL=��v��ʼX��@p{"�RC
���'�o5�~S��̓?`����H���e� �R�{�Klk���&2�O�����'`����X�.w�������~�8a��<p׎���Q�O��M�����%����W�t��R�	�
oH�i#қ�k�:�Ϳ��FJ�ܫ4��qe^i	`��6�����`̥��?O����.B�bܗ�L0ġ���&��:�N壈A������m׮����y�N'��+�� ӳ���m����2�����/D����Z�	u=P�p&FW�7R`P*xU����(I�6�❪�P�gbh�^U���+җĚ z1�@�34-iN_�6D ��`��yB��ް5�>V�؏��hÄ�s峲} a�<}$�!�D� ]bI�Z�(ٴ����rb��t��`��_���+F�{;�l��a�$����?���1�J��ig�1��ؕ�
��+�[zR��	��ņ��2M�f�_�����|�;\&7K��0�;#x�˴�F���������`�[�at��kuC02u_���ͅ���jQJ��lCuϣc�}d��-�x��K�r�4zs�����΢4+~q�?,���2l����H>���e��W�0������}�)���&َ�f�2�[��$��v�`g}�QpQTb��Ss�׈���t���D�R�FRZt�o�#�2z%��R�Ã�\��K�̸��#U�xg�������<#R�-�?E�R��������y=��(r���+���@�yE�y�����@S���i���^��!cVy�� ��%���
�V����UO��6�PG�����8�o�a��A
L|�T�Ϋ��v���o.$Ytب��"��a߻GNgE�g�|���{�����m].�l���O��+ˈ���!�"��x��vy�O)���c�c(}FO	�g׆�u�3aq9o�	��`Ui�	�V���^��yXa�G�+^���6A�LG�E��cO[�ps�P�/`b��^��3-�o�\C4s��Dv
�� ��,o��5[捸�^�ǁ�43�\��#��73���'��d� �2ǎC2�2���B�# �I,H��j4<���WK;�x�ϥ釡)����V]���Kͪ�6�4�Z�`��
3�I	q ��/0��N����kG��@�������������	,9�@w15����?��������~  ����P���J�+�G�G�9�>���O�?
�ڍ_���l�ֿ�n11{L��g�=��E���Gkl �G��f,�*i�ZO�V8���P���w�4 :j���P�/�y\+!��Qi�Nٳnz��N�<ݲ��;��ݷ%���5W]�_�Y�;(��ev��is5��N�~�๠}�P��`��r��܄����@Y��j�_frzѼ9��s��3cV�#2.�8����+�h�u�^�$�ϔ��^ԏW�>Sx�qI#�	i�p����7��\ξz��i�;ƌI���٫v��\��h|*Q�ʋ�^Mވ����AuPF��9�M��⦮��q�l����hBGAX��0�|h˛и@�	�l%,����B?ף�|���~f��}��1�o�"օ�YhW�Ȓ>F��\Ӟ�[��e3�e�� ,�#�
A�U�"��c&�]����K+��4�6�I;W#�2�v��T��-�e>�^�\&?l^L�P@[������PKb��R��פ6���.xB���z�6�cDa��9��7K�R��C.u����D����s��+Y��{�l��sh	v��N��l���1�(�!��6������懳/�Z�ۭg�Yg�Kv�V�r��^>aQ�S�5��\���(���o�5BO%iwP�LV�b���?�S��]v��:��"�\sh�T���F�P���]��P�i2D�ʮ��~�tR7Kg���l~~�gR&��`���9�=M!W�����FA�t%;3����J0� *t�����*ߗ�jr�|h"3!�S�#X?| �T>%<0���K���7�\"���Y߶F>R����BS�F.�Xy/\2�1U�KC#�B��CG�\P��N�z�*�n����X���6&�+MC�N[�~e�9��j�XR��d�.���X������`;q�:�EV�Ȁ5�Ub%�uM%Y�m��I}��F{TzT�\���e��+�8�-6�X#����n�ܜ��n`�h2h?��2�4�8i��ۛ�(5�P��=��*�y���W8��E�K݋z#��ya~ɕC�s�׊U@��̄t_��bb tҔ�H&�V��7A� RQ �ڌ�XmA�*��h� �;\C��e���^��X/�Μ��}ڗ{=o�`����h[��;�RΦr��kH7�m�{��S��l���2|���(w̾/��X�"�s�\*���'��&�%�,��ж�H˯9o4��u�g�۝�n|�A8�/J'	���C�������'�nr���CO&:�<n�)�柚�v�ֱʱ% �UQj�>Q�[�P�2�-�c���jz�Se�~�鶋��R!�/O�6!w�[����ZM�z/�������3�(ˠ���8�lH�.��ޝV���p�k3��������Ǐë��I(�4����)���E5��{��iSG>�+�9��2��a�#�d���D�"��ʨ׋xk*�C�N�X���M�1/�Y�6�};�'��M(���l��ͷ��Q>�Bޮ�	@��\&����O��Rs�k�ꅊ�)�*� ��
�mbN�T���_#tT%Ui�w	`.h�c65vH&ğtj1������Y��+U��l?��M�ȭ�I�ap���Vo�>2G�*>p\r��cPޖ��"1,�nxK���$�aĥ�?�Z��D?T�;�fa	��L�|mI]<r��^=�F��ǦdUO}:�픜��M� ��g<�i���n��^�]��S���l���������XQɻy������ħ�
Ňx;m���-s���
S��B�-"Ͻ�p�ka�?���0��nMd��
���x��0���X���[}W��0I="���-`Y�����t��H��y�br�JqD��+A���O��ە��������uc@��hۡW���嚞�����n U���c�𲧞��f&��b`Z�@��61������MIj���b5S�����pw)�J"N�?x0���I����)��PஓZ�#��|���������{xe1u�0l�xt��FL/�; �d���i$����nc�<���Լ�yP�pP����+s�?���P7�Sg�g�s�P���{�y8�Q4ۛ����@J����o�������ݬO��.�b����+4�Xh��f-��p���Te�N#]�c��A�]�:ʰ��`�퐯�x����TXg�9Ff6��~~uEș���K�<����;~^MR0
��oʎ�K����sU(�=�X�%�9�p��zW�>ZM�8�Q*(�F��U�^��m	�S�o4-��8�x�P`�W�\|�=��%��8cz�d���AZ*MF}y�3[bU�h�*H��_�6�sU7O̕胿�N��6�����ܯ ��"�k��Z���א�4�Q� �	b"��e!'_~�[������EF��ғ�v+UA��0��#��15�!$M��Է7�{ډ�"�#׍�aX�~��aO	���m�\�N�*�f�"GvIB���R�WIm�Ë�Hs��k�{��g'���t��������h���?�m[��<��5*�1����5I�EQ��˭uX#��sR��"���J�\.N�j�%GK۵���$�FB����:�R y>h��O��&p��� �2�ZRL��y[��m���'R8 ��?�w~��e\���$6뀎�P��K�qʩ�v�U/^3�vr���F��n�5L�~4��Ӭ���ɑ1MZO�v���qf\=M�[��e�KKc�!{�ti��Zv&�<w�m�v�4�1f��_�~@��Ѡ�@D��דc��*���C�!N̊7�$���z��?��؍�����V��hl�̩�][\QG&��jӰΗY�N9���%���tl��d������	��d�z��4+Q�2㮌�w߫�K6��;P�����Hcv��TtZtu�]׺�y0�d^YQbn���8�m���ǡڙ�6��ʙŢ�i�t��z�<N��n#�m�qgBx�_��]�,`�@)sdud];���j�����b�0�� q��CȨn��`�Aty��
n�� fz$�>.�b��]#P��ʼy<`{�Oqē'��X�%8PoXX��[�� �E�kJƥ=���n"Y�3�	���5��+�Y���,G�д`��Qp;�s�+��*��G��J!|΃�\Vֿ<�Ln�q�k�O� s�I͕^��:���<���0ٵ\�����1��O�bB�el���(rZ0g��jdШ!!�4�׳�"-H��L�H�br����8��`� ��>x�<r��Y�d�q��rQGQGWv;��½���2s�0�O7=��q��Em�f(��c���gN�0��Lwn����j��� ���xB�p ��+kNd���g�$epM��H�x=3s�Bf��$hL�q0� �C�@��<F'�{0�_�F̀d&i7h���x��[�f=��8L���6��T��՜�	�o�`w�:�t/n���Ȭ?���ߡ�l��qP���P�T�NvT���������Ĥ� ���XlxVHYEB    fa00    1d20(9ͥ`�|,���nӑ��z�At���_U6��j�)
{_�4�1�%_�dg�=�<�rlI�n��̇b �4xr��~ivΨ�%��{�"+w�3������S����F`�~Ir`�'���U�uYfd�ƜĈ�����؇�rߡ�4��̂b^���&J���|5ӊE~K4����DH�S�Q<��w�p%Uϩ$PZ�K��*�F�Rňbr���Tx�Z&J��~��ݭ���n�,��hF@���/�$�*�.UGÿ�0���	�p�
��)���(x�x�eH�D�zBW�xր;��W��D/\����r\�~l2���O�_=�%��HL��{�[��6��-ʠ{xh��1[��l�&؜����ڐ�*�Q=#�ۢ@͜�?�Q�ܼG.'����1ڵ@�@��Q?H�dD��ݶ{BVAi�V��8qm N-��T@�.5Ɏ6p�Ɛbǜu⳱�����ў���NLT�:���i�y�I߰1}�ǳ�V�������eXٌ��k����6�F�E�������!��(���a�`l��:����4��/�p�	�����8�|�#I6�P�[+P�꥗�~���.&N���)\��=����B�81W<i�
�)[������Q��k�#	5{}�Ѩ	�j�㵪�lH=���N�d����!D�aM��q�S&�-5�����8���'�rM!˥L۟+�,��M��A�ہ���)�Ŝ��B,D �]��h�,���8=���B��U,Z�g@V� D�s�7JlVO���� s_�l�B�z4ތ0)��P���p�o�� 5�� v�<c�U$"����2�I;qp�k���r��S����L5��O��T����������Vp[�k�CIjT�-D���F* �!-Qu����J�Ot$�a��{�z%nN�\�"|j��g�x��E�V��Ss���Õ��|A���`���>�ԫ:}��W�%je��{u�a � ��Z����H�]�Wp�@��'d�7Wۄ���|�L �`��1�|�[ìz���RΌ8�:�%��+�/�6��Ԧ�_5�v)+�����mǑ�wG*1B�h3Oyd�b2����C@����^�C>J� ֍�G�-�uF����~<�G�-9/��7{�R��l*?��t��:����2��H�Lx��~�1��9����2���
^~���f�z�cRb=�Gt����T�x6����)Ҧ"y=�F��s=*��l}7^���h�H�6������T��sb�TY�'��]5��-O��m�Ps�|�����r��G{�Q-�(.����gc�T2��[�̔V��w$\bV�B�`�� E���?�H��A��2Zʚ�o��J�N� �;.�	#y2������ʧ`��1�Q��,]��y9� ")p�bs�$��K����h��/e��U��?�M�D�B�����@��2U_�@Of��ո0ؒ/��C%�fB��5s�+��hzTE^Fz׻���C���ܬ��YI�����}+)���KӬ����-Ì,�Η�a?�m~�r��a��.��W�U��q���7$��*�Ƙ��	J��8�d�0b�_�IߝS9�H�Sn�׎�v���G5��ќr�D#sV�e���|���l�-�BP��w��j}�=AI<o��J�x�1N>a8���6îXDM�uh҈�/j�%��jE��9βq�iH�ȍW�mY G��<��N3�)<����6� ��{���f��b�^�
��=>��>$%��j�U���������Q���ʁ��V��H����T%
͐���j���'tk�Kd�%�VS;s�����.��qI�c�\�LR�*ѕ��8:�����[?��wE� V�#c�O��!�%X9����F|���q�kԾ��Lg��#cYCT��𜸈��}y���Ǒe��я�\��3r���4��!.���YJ
O�;�1�@3s����h��� A�5��yb��S)��-}��d���n
�3�'��V7N�,#xEU�������Si�¥K%y��m�(��_Zr�:é��C�}PdX�]�v�#_=�E���ʕ�����XU���Ȋ+",��}ieCko���Ig��'���;��eDL�G�ъKv��8�$��bs+��͖$���D�JO���]�������kA6h{�vH�MFi��Wm�@����J�^`�6���zމ���:�o_�l�nЇ$��q����j) Z�*a${Q ���D�������97w�0"[�b|�}uYd<f�o^���MVSl�uK�V&�6���5XT�]�*&�sdTNx�+V�1S�6�"�OQ/�*_�u|�D��ElA(�;����((w���	���4G��Շ�Y�D���qhzk�/B�o�˲I�4f�>o^���j�{W�C�w���C���e|��	��2&�	S �F�s�:�?�����JH �S��թ�푆��
�m˭_!������P5ƃ�m��W=�榺�5�N}/%1�=�-O��	����6&����Z�7���4�m�ڥ���%��w(���MhĂŇ�=M��W1��غ�,��r��8�L:�Sq\7�l�)��x���<6e+0�d��~���Д�,XKX�7��?�4��T�@y�����:�<���nK��w���"5y��O��L�BS�Uh�`����X�3cgY�m�'����&������v��s[��*frkA,��x����%�S�]R�j����!�2�8��|� ����\:4>�
��?�xA���Q�4��YQ 1jk��-W7���C{Z�땭@�@ ������������GK�w]Ř?�h���v�����C���A��6g
�^yƔ�gv�.��y�k�ZZ���PE����$�)d�5'��ři�UĘ\<�Cن8\��ݸM��߽KJ�Nb�8 6IO�6{�f�Wĩ4<��ﴕ�in�X/�nf�P��3/.�7�bߑ�x:ز;�y�+���"AE|�2mrз������#�ϙ�ތ�㲆sՈ S_o�[zt2:�Zy����A���r��C[��v�4k*���=�qR��v��;*m��6I#��c �m]�����%���Ub1�o8��}5��C������ը���!6L�.���WMpS����/����|���_BJ�ár�(����_	B]�O	7�*��K�!l���i�ln* @���tJ��]�D%�|U�g#��z&��⵩e��M��g0�m��[2�����2,�DiՔ�-��� �����ZP/��)�Ewy�t2�O�;���Y7�TL�ô��]t�6kpKD�{q��L���G�_G�,�dE�>9ܬO�#�,%��Q;��r��L�ir�,������iF�2�>��?6�xu���N?�͝ߢ(��2)�Pd�td_�[9�|�G3�<�Q��Ӳ�llXm��ۙ?���fW
�X^f��QI���@d�~����l�a|�
C�j�9|������;�3Dr����򸁉���JY��}�'h��D��Ό� ��5m��>�}��Y�󆒍��C�9ۮycp���!���K��N��ۭ�W��I˺N�k���z<z�w?\HI�u��».�Ύ����s�t��J�^P������������A��֙����q ���VVS׭���A�T4H�D�;#i��9}�FO5W1}�����u�p�R�c�� ��Q���|����^����w����U��f�#�wVpvSpʨ�_+4q���Q�랸-�c�/c5H�+^\d���f�R}�LM�2C�5�S���:������G���YR�gV����c�.�|�{�T��K��3�g��2�b���@q�	Y{kGE�-d48�摹&�lcDO	��Ș�?k����f*����K�ix\F�|g!3�C��MQ9c�a_�L˪�B�s��X`O������{qy��}\�?������ZͱD��Fo��Y����E�.�"�G�
�J����Z)悘zГ�� ޣ���F)���z���W���X	�T>/��غ��k�H���7���l��c�ǳ��f�n�쀟���@׳��%Z���%+;�� -�;���I�j�-�ݔ�����9���*������Z��V-�Y@�.�v��>��,�|�q��c�~�-
���A"��z�"q���0��n(��K��W����0�I��Uq�	�ۧ6r��r�GG�`�ܥb��v�P�uU�����,�HA���<r����l��9z�B^fŚ՚s�:��*:������Л46 B��e�Sz��/fK���?��P�m��Se<h�(1�K� �nk9���P)�)�U��G�
��<�旽)'8Pr��˲�p�󍺸jV�;�uq�ZW��[Z��O̸���"�-T��v�o�%3d�	����U����`C��	|/��$����ՑH�p!!A�m�/xidh`��U����kB�#Ҏ3�MwSQ�p6Xfim�䲚Qn�h����P�G��'��Iq]�b8���_����m�������ɘ=3��C�qf"c�8�����`�ȩ�eƢ������\Õ�\ku�-�nG�#}�YE���7�{]�L��vD��OA����,.�C��U4�ˮЕҿ����D���z��+h�Y/���Y�!�R��\J"�=%6��A��UI�57S�EI��-1��)�`#��'�4XOX����Nk7�.��Q��8؂BD��J�U{����I���')EK���������ŵ�5	�ʻh1�?b���j�I�,������i�JxX��3?G{1��_s�y��5�$�}͕�ˌB\�ZN���"<��َ�`�'�Ft
������'���D�R[�$NW�� 9ǈ^%j)�{��!�!�r�8S�]�fq[�(~2� .�Z�ܪ�xD�ei�<m������^����8��3W��I����?$Gt��'O�[ڎ|	�w��� Y+�J������5Ȑ��=i9k�J�Ղ��O�?��ʥ(Cz�7s_�%�Э����1��Q,y|+-!�ol��<=���ȭ���������k�B��.�R����a��A�o�Dú퇖}�g��h6�*%��%u
�"XG#�x�D�?R�~iq����D��j�d?�e��{L��k��%�\ ;�o�h"9�`���+��e�:��9����:3;��_��T��T���9)k,�WmG.������-"3���T[Gn�%j��_Q���C��14~��b�����S�.D�����}�w2�Nᾴ���P��p1��̯̖���ܤ��Ρ�x�{��t�`�8ͱ�sٵ����Z�.���� IX ��2����w��G"�t�1%�Qv��zn�3ʬ���PC��Piķ�\�/�m������NKG;4�? �r�461�	��f%?���Jv�}Z�*�IB?zd6�0"�o��r����0�o������Z���6�b�����0�eɑ��Z��GQj�OϾڷ�{��6���M���b��E-��~7��
tuJQ�]4��#��է��M95��?�#��p�@���}��7()X�X# X��$U��7�z�%�̶_P���X>�a�;}I����a1��f���m-��ϰ�Ϧ�9��G�R���IP��%��
���ub
~���#A|���N��dr�E�]<�[���I �Y�<��?-Q�C#;�޿3�nx���&��B��4W5����hC���>�͑_S������򐈬E���\ǟO:�]Q���h>��|���ݑ�(^E4!��e������o&�P�9v�O[�7��0r-�qŤ�Ko�0��ϟ��3#��*@��cChƍ7EbF�3�Ʒ�lur�J�Yt�r� c�Ƌ���!�T�?��n�#��^��=AE�q�vF�q�̉���t�/������Nu�y��`�$F�Z�T�tX��'6�[,�w������q��Z�� �����(�u0})5zz�*`�}�Ė��B���q�y�oÚ䨉�A��7����f�_�k�2�+����`iWP ���Y�DS�
���k��Lr48a���դܨpS��
?W�������+��W���v���,�JF��n-{�\�i�sÞ�x���/實�	�� ��g�����0���&Ƴ86��x8*'-| &�����I���0�����#���r*g	�^ ���█��O]�10�_�A� ��� ��L�3B�~���՗���Q����8"cSĘe�hSFԲC��*�x�6q�C�C�Sn�-]�?*B�S$�LlK����w=�o� ���J���q�����"ۮ���(�:;,<voظ�V�vM�&�L��fX�P"��y��}�o�X~�7�LI�)L]�$����q�>�O�� t؈����뾼�P�����O^�sfe7{���G�avKU���:���x	��H��ҹ\��k�^��J� o�!�U8%�h��W�� ����'�9�)�P� {w��#���X��kV�}Q!Q"�{��5���#����ͺo���h� $v�4��c;�L�IZ��O��z�=C1��a�襮�D+NJ�ak�HW%��j�P.� ���靹� T�yOCVC^Q`Jy�[��i �d�\)�����n@�����n����8��|��`��C:1�CC�(�u��C�$�㵦n�*� ���,��4��Ȱ-�������_�� ���#~������������A�l����t}�J ���&Bx���#�>�v��y�΋�8��?�,�!�ʞZ�_{X��
Q���n�F�0��2qخ$8͙A����%8[�I�L�^͡椷�j0xW0x��b��_|,�h����_e�E���Gs���*&c^V�D�`Y��t�̞~p�r3�P"u�O�^ȼ0�	����D�K ���h�ai���<���u�eQQ��j���i>Y1@�)�!G��ӲF�h{1$�y��1w���^�ܵ��/n.��۩��t�Ck���*nA���
������bş�M�8����j���)W��lOx�I/O���Y���!����[�m/�d�-}n��(��ͶX3]c�/]i�IH5�ܛ�ݵY,���^�RZ)v�7��b��=�Vg��6�H�JLd�!�J�fN�B�&�d��B q 1�ԭ响۞K?��g���uDPS1�r4��<d�#���q}c��>����%��>����S�w�(�8a)u�ǿt���P�m^=N2Ɲ^��jkQ�C��ͅL�20c��7�Sͮ\%p̎��j�{⥉Oh�P��T��_>Ȃ�ʗ���_��W��_�(�/�Tm�
�&����7t�[*�ॳ�XlxVHYEB    fa00    1e20iW'9�W`��e��USY�����|��㴹�l����ީ�H�Y�D��9	}K�?���
D{a���gK_o�Xk(��[�l�O�ѓ+��f�褐D�mbVL��a�+�
(��a�w��h-�>�Z &�S��J^��%p4Z�)�e�H;V�=*2o&�F���"��4�{�4�Y��ѣ�eՅD�l]�»��l:����p�)���)�#Ay��x2g��/�N��;i&Z���8�:���]���W�xs�r[n ����[������'|76��	��������V��ˬa�O={ʉC}W�}�Mv[�5�i�|�Qt�Ų�h,	���K&M���(��u ˱�|���`��},ufv��Gk�=�m|X"f�#�0N���rq8�(��4x��:V������<$�htp��.���+fSg\C&�<�MQã�8g�Z��T�Yvx��e�X�{����z"HI�����m�v��*F�s�r�����Q�'x�y.&���@q�v�K��vq���f�G���=Qa��)�@)�p��1�׺��X;��4i�H�AčO����]~yу�z�(:V�ˏx�c�#�V���Iǌ���2J��I}�_�6�E�NtNl��@,�L��W�����'�R\2hI�)b�FsE�7D"���d��EV����0ْ%�Е�xvc
���f�>E��Aīgp>�{5���w�����ݷ?�[�:���ѽϮj!VB#l/gJ�>��y�����F�������%ͼ���=���t��B P�]�_D�JrM���~��c�����2�$�R�e��:Huuw�N���Wrx�����\�;�0���o�}�VZ���}��_��U�Yϧ�`1�#�̉�+m��7�tZ}o^�n�jTq#��/8��>N�D�ډr�X��O��	s�9wM���|rkt5�Y
��Ee�X?���<��,�e��I镝�i��Y�BPp�}}��.�L\��i�˰��g��]ʏV.ۇ`r;A��y�{S�!(�< ,b�3W�)�vV��=��%�b�C����C�tE�/�$�veGl��7+7E�����j(��#w�s5���*�������R�y���(�8�,�`sE�~�D����b���g�Y��y��t�����l�U���l߲M��8���6�Hgy�I�/X�[���nW�b�|�a֜@-K��*s�l͉o�Ș�SM�*�߮���O4l�M��}�!woU��b���q��2���_������
��뇴�ՊBJQ�cpQ��7������n��w�l��+�}͗}�JE���*Tx�>�����8�JYY�8#ܢ�n:����;��LK�FQ�?�y���Ԓ~@ɥ�����`�[
����5+,R����*M�#p#��gqW�x����h�J"|�/d���L��[��kZL�j�-��%d�b�a�@jV´�1Z$U5!��8�������y�p�Y���3o�Fi.'�#��$��p�M���x�Or��Br�5�γ��W�<J���S&����GP�YE�n�(��5H̒�-q �f��S�i���VL/_�\`�JYȲ�j�t�H���P�<c�|���D��ߑ�s������e�^�7�$�r���sFq�����mu��PT%q�5�3��>k�gs��0� �~��2���Z��x�rq��h[����D����������A(vs9< ���΀��g 僼j4��-��:9A�-
������僸�&�zq��ĀE:Zŵ�V_�&�tq�ho�Dh�\�fN��l�A^Qd�=?m��H��B�8��wm�>Z�͐q����)�6�<�_|"�CF�#������g�4�2����	��_��
G��/��_M.T�w�K����m-�3D��Fη��~��N���m�FBw�� �5��XU�H�/h�w�T}5��	A��r$a�g��[�;Y#)��m�sa��)<�;DH��XtVl��{��U�X�N
 Ʋ~/���"��}��?ɢ�t�toqѮ��HƏH2z�AW�s�$�+C�ܚw�̾�#-�(��2V��}>�y��,q� ^�%fJJ��v�e�a�X�yRA{}�zy�;gv����µ��#�����-fT
�J�\����b}�o!E�[��@��12[#��|�����͆T1�q������v\#����PO�w�o���I�q�%�׋R�N̈́㷥�(���C���!UI�r��}�iM��d��F���φJ�Y����3\S�܉?*�X�E¹�I�@�4����i�r}��#(Q����M�p�D.�)S�VׅG�(��O�F��L?��q�7�<�FՋ<оh}�v��k����
��>4G� ��[WÔ�_�o��o����2���ω_h{di��]��3�<�d�qx���gh�ӁYG�oY�ԃ"�И�Qc<��ޓߩ�[Uć�B�!
_���t7BO�s|�[�a�XiT�¥8���@��D�-z��@��Õ�{�v�.Z��oH*ק�Y�L²�P8�&�����A��|��V�a�� �da���b�}�B���]��z�wN�M�);�=��a[�t[��\�3�f�.����o1�zt̹L�"������o���)~��q��j�����F�匁��+�&a(&��l�d��8Y�x1N>cKW��`�N(htW�)�f��<��ݒ��Lk�~_B�;��Ґ��m�G0>�ԥ+_i@�� �0�^�"�nO�uP
@9�A�x�b0>��Gd&��]E�c�2�m#0���!)���*Bu���9�rײ�d�
�e�qc�	k�<�%�e����U\Cv���I��2�oz;%����"����\$U@�[�s�ܺ�'��@�������}cx遻�f��W����&��7BM�}|����(aFZ]�v,E͈UOr���8|��y�r�A|����U�^%��l�L:#�0�>�r��P�JYI�
s��f�&��Zx!N(�蘡ey��5�1N/,?�IGg0m�F�5��P1$����c�x�)��^��g�~�}P��w�/���� � �O=�0 �Շ�i,��kV�7<G���`�sHL���3>99IxК��u�ʖ���p؋n�j+4��.��g���:��L�����`Eo�4������Z/w������v���)������Dd?NU�\�իYLa*�@���n������E7]S�U��=�0;�!m���ߎ�q26�g���C)B;r�G��|�7�����ɝ}W��-�YG�ӝg�51��$@��}CrgCcs+����豠HZ���:�<���b�����$-�Tt.�S�c�����x�-�~���OBY �a��
��v�W�� M�'�$����^�'!;$e߄c9�c���e�"��ஷEHz�lhÒ�=�ls�G�
T��4���_������t�[�Ob���������3y��k���SP$LS�ked��_���F-�I�Ha���$\���>̎1�01�%��Sp���c=��*��"H�5��y����T��'�m�82(Ճˀ�#������&C����[!n�a����K+�y2c�WG�^ɧ��% �晶@�T��L�zC��2�f�	���%P\gˡޙ����2��_1Y������l�٦��$���`��X#���@��9�qֲm�w�M5?��pi�/�N�u��|���9=f�4p�|��w�
%ȃ�wh�j�1_�ю�X�Hzp4�}n%�4�\0�v('���f�2.�� زF�\g�̓�K�W���g��v�R�g:'(�
�؝yv�s��9n��V@����m"��X,u� �p�1@9�<�k7	y\�V5/-眹#*�^����.F���̀�L�����a���	�O�]/��S��W�{'�c��>�h{LۭZg�IÚ�¡7X����2��kǀ
�4.T�.k�p+D��;:6H�QAr��Z�X]�1iv7�K+�	w�udd�N+"�ư�(���щ&B�(lu��ñH�N[�����g_�� ���5e}d�D�OF� ���Ps|�w�]6���@%[-a�6����?����Tg�+�<�Z�<-�"ܫ��3�.��$�����G�n�}+��g�6I��-�����}�>ެٟ����b��dO�H��C!���#�-`��<JStMpR�4�#� Ot�G�p��!ƒ���EX�D'e��p��+#[#1Ne�����j�NV��[��+7�����WU�U[��9.����O5�6���C�Ӓ.�8�0b�?�@��j��a&55�Ym>��3c�o��ȶc�q��	ܩ9��	��z,�x��A����͗w��u�١��.d "��I�"]3o�l��39T����nT�s?O�,���} N�E?�j��(/%i���� ,}S�H�N0���aOm�f�\�J:��H2�><����o� �hq�i�V�	�S�΢�Q�T���w͐G���f4��[�&���3\��4/��.U�ڨ�����γ_F1�'ے�Ά���6��\�a�)7�$�6:���x�	���ʗ=��B�lF�q���s2N�����D��ީ1y<��L�D��gb~�X4, �}r��*�m�s� �C�9X�b���`s�K����Q���d�'�Ss1��ӗ�����7�m�SƆ=�����[����BI��%��`w���.N��d{�^L۾v@�οeo�y�v�r؊���f'��`
��;WH��6��G?:�/O��q�ِ���G���� 饢��c��=��=����"�Ѳ"��p)Bcb�9>�ziS���K����	5fКĦ7��lt����[+����f���t"���$Cק&u���h�p�PM��t��>+k	�O��)�^bK ��l+��֬E�N�m�Ɲ�k'��cO�������d������M�%��wJ�|�l,���V�*q��'�}x4�"��.A�^w��fO꿕���7�Ҋ�c��MZ�Y�v���P�G� �߂���^���uR����61^����PZ������Q���/��4�_�H$��g7d��Ѽ��k�i����[�e��pr����0�9��8"��P�zse�*��T��qdS�5
"\՚/6j�.�����|I�ӝM��6Vs�;ct����R~%��h@N�Iqu� n_ꛝ�l�����N88��t������r�3�*���j�o*������cp�r;��5�ꇶ��䩞F�d�ʔ�&���Y�>Gw�&yB�EtQ������q_i���\T�d�&�]#������K���畝����P/�߂)�f���s���{&�,�I�S���㔠�J�+�%]z��4���A���� Q�~�r-_#g`��Y�בM�(�3�b*@��|VR�%`7�MT�T��(u%�#3�4�%��KѦ�S̳�15��l�a�		s�H�V���oAab ��X���ŇIB@"?��g�����F>�x	|�5�8v�sY��^�+�l,p�`������5���A��3�����k�������C58D��}�4�3�Ė�5P���WQ����Gº�T3W7J;��ۙK&ѐW��bd���aq��SAf���\���8-���Y%��k��>��󠔠D��Q�hz[�ۿ���d���^�1s[�2�� Ҟw��>S�V@�J��s���~ޚh�MK���B$�t�N��Hj����Q����!�I�զ�c�El���5�$�g"g4�A3jѥ�^�� ����V#��u�{XwB��#΄�1c�z!��z�3U"E*΁��Ve��9	OP�k�H+�8�l	���+��rohO_*�:��mݣ��>F�+I�,�/�(�ɣY�&�|������������/<�?���#rtT���ˇ���xC���^�Hq������W��L(�:��~�]qW��v��!n���l�����G�� ���Ӳ�Ͱ�%��$?�y��?��~Z�Z�%Po��Z��˄V�.oxZ�TH��<�:�s�Fg����
h8TY�]��)6��g�a
y�.:�ʮ��g�rT2�ء�_S���ϣ��T0��#�d�2"nk�Ěڳ<�#Hn�h�ʊN`pz���˗���[��RЭ�&J��Inq�!�ۣ�`C��m#FM�e%hZ��jPN-��B�e�������m�H���52��t���N㋵�Y|����^�o��iڜV1���z'x[��ؐP��)\�Č�d��[��ˌ�[T����,���@�[��G��U���(VC��i�f�ﯓ���לI�V��e%�i�S��j�%�=��IQ�q�\Y$N���2��e�گ�l�bY�_n���$�t�Ke[�g��]��hM�UO�+ଅ����w��|��d��/�-����b`�v�W��"M� y���0���+/�3�/��7Δ~�A�73sx6!�Ӎ�j�i <|R�<P�X�E��E
���	W����}Z�ġEf���-�1ϊ�F�+��& FW�(�����A�w��}/���:��뙀'���0nO�4�շ���'�����O��6��a�,.�� 렺ӻ������s.c�ZlVՀf�MI�*Fs?��aӽVȭ8�gOtߕQU�!�R����L�քu|���m�l �K��6~1����ɛ�8$6��b�8�а�mؚ>f��(�@�6���O�(���K����mY�e P���ZN�߻�cI�>���	�M57}	�c�z�I��?��P"���{6u1��e��&.�P��F��ج+}�9;���]�9��m� /�T���ԅ��Ԫ ���xЦF����l O�}Ik�8[�U9��qz�n��k���o4�.µ��~��2�E�U�o��[u��9���8?+j:u��(,Xs,�����4mB�c���QJ�wVUx;~�;�+z[���,*@�<,o�@���c�Z�|�qq���i�q���X���mna<R�&���C:4�
�/����1ͣ~����u��j%��V3_��e��P���#gB5�֚B�4��#�@E�5�$0�Q׋��O%u����d>���wæ/�$YT�Q+3"��GJ�=���2Nx~�*�;`P�k�ݨ�����@�CH�L�M���z�a��,�����T��`[[ċ9����1�����3'��WJְ<��h\�u9���X{�ն{�:v�Eqw_��
���!�D桉"=m��º����A�#��>}��}�fq4I|�Ar_U ����O�gQ��GX?�xC����sD��k�ٕ�A�Hl
SW��!�	/&��Ϙ�(Rv��s`��̉3RX�C�h������܏_D��yԝ�	�)�
,�N�(iG�N����H��r�Q�AT�x�}�
A
V�S�7��U�ە
��ʭq��5�}9{@T_���No-(�釜����G���v�69Z�j�]�4�]�(���.j�gh�e>��8�E��B..�ceR�f��#�
�{�oL����`�C;	�?���F�ŋSYu�t�SS1����S�0��^[g~d���G�<��XlxVHYEB    fa00    1e50���O`r���R��w7�f_�ZL�
�`A��H�� jJ$��(��3_��Y;g�$F�ֺ�z�DN�	������� I\\}��(^FAK|Y=
�r.q���Mc��+D�r��{&���ʻ1�ĳN����f�`�8�s�=:�;���ᆼl�(Nm)�3�:��2�Q�ܙB~!�*�;��<)�7�4��f�܏ U�/'(����<�_-A. �p���D�y@Wi]�h�dc�< ��O�_S�u����V����|�*����2�&[���7
����X��o��R�u
!t���������� ���T��ծn��?3L�ݲ@\
�ˌ�%7�d�xj��������Dfi=�M:bT=qx.�N�ru���2�;�J���1�͢�د����v!�,o.���[}�K2L3����+g=��7�F���E.A��g��js���:����l^#�K��W{64�]+	���*�H?f�9��Ǉ/.��
H�-唞����+]�@��BI_ݓ�"�������R��#ZJ�d�.G�w�$��=K�B$����.�ߊqA�)Eb&�ƠT)15')�s�t!5/纋W��s�uʔQ��`� ��v��� �i��K:9�ai{R��=���^E|�ܹ,k��EQ:��&�*�'!!����}Y�<T~���r�U5���w��H�c6{x ��A��ua��䳧�<;���PG�w��/��e�8�p�T�E�ݍ��V�&���f�ũG�R ���^�Oz��Ta؃((K�T�Ĭ�I���J%���A�0�1�8�JjAbRɖ��cB=�<�0���s�F,�έ�����W��M_Y���J��G���06� �u>��-�6���X�M%C�������Na���j���X�K�	ec���;�N�K�O,x�x����*F&�IY��Y�qǎ�X-u��*�k6�g���$�y�CzF�^s�#�|�t�B����6�+}�=�l��0������D<ץ�f?,H^��퇪�JDR���@�%��q	�̓+��A���ڣގ�$5�%����M�Jy���"���=�����}�
%�7�v�2ykG=�{
$$K^�Ne(��d[�A�lOvg��5n%�6�~"Wh���"�z�Mb�Ũ3��/X��q��M��8)�i��I��*kVr�ᫀ��z��lQC����X��aҲ�!�r��h�.O͈.|���sb?���E�D�:O���L&gt��������"�"�8�{���7������� �&$�V����6:�kU�q��d���z��W��1ǖ�ŝ����+h�x�1H�2X��6�Yݍ![��*�]����3N.���ċ>��QXq�p�}J����:�����������"/.�Fx8��[�"���z���jwğ�	�5JH���#��;�45���w}hjU{����x�ѧ[�"����<=,%�╒$ �w�;hI��Mq�L��qf]G�f��O�7?Ir����}9X_�-���;6� �R��a<��Z.�Uk&�#T���2r6�m8�Rody?���=$l����
'U�ܹܰ�O��3�vW�F��2r#Y-"v0��;K��!{��X���d\�up[<Cj>������dn��:�8�t�0Hbߐt-=��ƒސ��
+�뮡��C��G�!׊c���������1��HoPf�ł#�k�?B_$ǿ�ٹ�� 'HV��ˑ�v-0�0���-�%0���=����wAUQo����i��ݏ��lz�����^ ����-}z��:�ە�ˎ_H���x�~�|0��/'O?�� �0H�
%��e`�^�ѭտ0�J���Ǩ�rӈ�`y�(<��e��)d���x}�7k�����*��s�԰'�j��jǝ�s��ۇ� ��m:�3j,_��� D`��c�ZRy�����eNӒaj�O4��#��(!j������1�E��.b�r���u��8hb�ڕʬlķ٤�Z�3�v�p ����5n���P�ۥ������<���#�����lh�צn����s*��=����S)|�yy8ovΟA� ��f)��}�?�tlX�,[�xtr!r�)�Ek�=�<��A�(�9� �{�� %���g�����-�s���%q:�\�nR%����uk��t4��-���9��i�G3����1�W�}�vF���n�c�b䁚\�7m~9x��U!ߞb�ц=��؎���*��پ�m��X�c�Y9�@al=�zC)�#R~�p�"�l�=�/�_(Jr��)�2�z�K=v���v������cm�fU�� K���$D��E"��!m����B&M���Wv
�9�j�͡L;7������v�$;1�;߉Uot�s�8�|�n�&��90����e�n�B�s���m��Y��/��|tl�t����6�ITqon���6j�4q�6~m	������,�F5%{��0�ﭼ(}���O�u��W��Ǣ�3�곟Q_Gg+=޶�]�x��Es���&�m�^��}B�4�n�۱�8}*<�l*�5��a�m�F�ˋ�a��G��a�������#kRm��+C��{�K�����]c��U�g� :=���D'ֻ�<j���	A1���N��"�lHx�k��9���A�}|�{oh�<u�grҙk5���/	���g)M�a������K��_X6�,~ܗ�H�:���*50�0$���<�s�Cاʩ���`*h�CY4��l9'�b����u��$�ŷ�-�m�x%6��Q�b�wr����v�ĉ�-�PB������t+�G�  ��'ZS"��B��*IZ�]�J�7��Q�0�zk�	��B���u�����F?�)�R�V�=��T7���`�����\Dd��7d&�"�X�
?\�0��j�o�1U�xV��X婭��Y{hd��<��`��B�su���g4y�ҋU+���)�Ϩ�p��i�V�����L�+7>hO�>�(��:� ��Ѹ�K�1$�ϿdU��qP�k*��=�H�V���a^>52�+�*�u�ho�)A;;�~B��{���Ra!'�/^"]�*��VEbO$�`��4�t*N�i{	I�6Y/y���{
�,�(����Ĥ�ф��P�P�����q:�#�8\+1�ъ�d��H�:���r!����=��S>O2?��)Y���Zh[��*�՞�ACŚ���"���!:��|�}|q�<b�/ �B�R��p��k;��_S�i�9�1�MTpxBp�+(���J���V#O�\�{��R�bg6��v��.����6���ܯ6��$��)�.ܶ��M|�Q�QG'��	J�O��m��]T��PN����׭l���Yɛ�e���v��v�i�v�h����v>xD>)��Z
��V��{aJ9J�rv����-��طӓS̱�h6[qpp}��f1\9��i���/�5�,�ݱOS[��"�ݰ����{���qm���:j^�$>X�(��u�Q��+�^��X
#�5�0����]�8٩������$_�v����(^�VN��K� )5�~m�;U��� �%d�\ר��\��!�ӑ�c�d~������6�L��[�|���Z`��9sX����U�<V�6�?f��a�
*a�i2%v��Y-�B��x�l5<	�t;܆�k{��x����h��\��D�{���|��������*^��uz�C@����~�f\a��l%�L�	�R0�|竴Ҷ���,W�U�h��zFO�U�C�ƪ�DUI𩷿�LLT���6�HTK'��R��|��M����>�g�1P�؟��40���)��4�}-��i.^btb�9� /�d���:�A�-�W9������L�W��(�p�C�B���(��^�~��O�y�"��qj����\:XQ͊�\����+a�S���|�e=�O���̢�}��N���7�:ڡ.���ai�R�mz�fi��1����� %LE
����n���Ix_u��t/j�?jk�dk��݊��XJ�:�=d:�a^�+�еu��@�閟����N r�^@l�}�$����D�8��B��c�����B������B��y�ݡ>3�a�C�R�'�Y�� �"������&m�Ĭw �6d��F���m�~c��g��CrҾ���s��.np�+��*]O�����cov�?��:I��| �(�b2�N{ə y����D�	j^��9|��͠?�	�j��ԁ�ٚ�r�0��4��� ��S�i�|mP���9!��%�-�F�,w����]�ڥ�����dOEKo3���Umh�)��鷫zdm?�_�#j^��IP��.[,x5�Rr�x�̫���l?S�ot+�{�`ie�>��p;����zvnd��*~��3�+4X�X��⢲�I�A?\+�t[��n+nC�����<X�|���о�qJ���?��� ƶ���ۆ�������M��3!!�sq����J�&9fQ6���p�g�-V�b��)��U`�j�Iʃs�ٽx|W�!_���I�mt�
M^�s�5�:��G@�c�S��Z�,�8���Y�M��6�Ǘp�Jmt��D>���̝iA�0�A*=M�2���Ӳ_��s2b�!��1%��3���eQ�<J�z�:�A�6E/��"�����d���c:7��C^i���$Ӻ��U�/��֧[RT)Rq��0@A�u.�u�A��"��������'��ضìW�ZJ]���se����{~!���H@O��]b��F��f��~�jf�� sHT3�@��[�Q�la#��	�
VRq�/b!M i*�Q�`Zɼf�'�x�b���*�g�w5��2��2��������IG{�AC�^�Njm���ދ���Y5���8��xI��%�5��'�r8Zh�/���s�<P�Qn�p4�J��[�8L�QT��5����-��;;��&��J'�[3hn�i�)��cʼJt�������l���z�^����gKp���d;l�:�����C�,�����&0�����j<�f��c;44���	h�td8�X�]:��~���fRV��ﶃ�g ��ƕ}E�q"�tY�yڳ���u��o�Kr]5������"��+�T�H[�\���? �<�2�S���2��0�����lmw�2�[kL}����:���B}��.G�`C�"@nS��-��'Q|�(x�4z���5׆��A�Z��i��ˏ;8f��ʟÀT;i�Q�%���V�d!#���XuK|��-L���U#`�J�~�|��� n3ȌP���Ж����
Y�}=:=Z&1�{�k�q�?���\KX*��< @�\A�=&���Q�X
ð�l�*u���� 5��'[U�'�z��O�٨x�ZK��g-4��o�:�=��1��D��΋���GQƄ�s�>���0_��?p��V������	�Ƶ^�Y��k��j?|S�2��֋�e����J�)�\<�Wy�QC��+�u�S��U��+J[�W�:�6�~տ�����8��V=��J�Ĉ�����	$�"ڨ�{�-���9-25x[���ͥ-��&�z�I�'u�H{�g��'K��d��Jb���������F+���D����1��Q��@�o�k�J�)@� e�s��{�������]�=�/H�nZ׊���5U:��tan��q8�%��`c�����k}�(S��Q`� �eP���QPN?D����j��oM��[UkngB�[khQ�P"u @�� Y�:œɅ{�:|[���\3�-�{#7���$t��T�Z��Xu�l���d��=�B������.z����G���~ ����VӬ���ւ+6�P�W����,8�ZrYF�G�B�j}U��<��E�
掝��1E������ ��BP��4�$� iR�]�	��kmA�� 
EF�|�%���h�5錴�dV�=���
�W�s����4��o�驾T�p�?f����"ʁ86�Y:�u&��L���<�K�G�1�lY���_W��)ɖ�*6Y����C��(���)+F*ge�a����:��G��.��f���6��{	���8H�-�h{�rȂ|-0U{���&nj���/b^��
���(�[&��ގ[+��_�`�҄=_���F�������z�jAbe:��Zi��DkV)���4�m���>L�������m�[�g�#�rF�t��GL�^�l�=	[E�51:�%G�nM}=��F}�O����1/��-¸z���IL�@�ٓ�Ѱ^��K<�,�kѽ�H�)�I��Z�"��gHb�d�{2gx#��$x~���
K'��ݰm1u�1�&�83�%�+��|�#1�W��"ֈ�XC���ʿ�ܺF���p^��ڴ2h��:В nz���t�?i��������⃶&׃u$Lp�VA�dL��V�"-?b2�z�����B|ax���V�0�h,���qK�����n��i3�6W�JW;%�������h��^l6�~�pT}7�|+7ۨk:�ĪJ�J�0��%�;�����%3��p9o�]�d���%t��g%�3���4����Ti'��*�wY���I�c�b���%���$$��/PȺA4lV�9_��~4ER,�IxI�EM��0?�K���<]+�00�(�7��1Li��>�%z��ٚ��o�Ie z:fF4[�3�B,�s% y!r6pvv�Q��q���0'
���<�����Y.��4c� 5�e��,}��.tl`M�m���";,�ő}>�Ʊ�i�i?�W�R�l%�4ۯ�ܒ7ID7��e��KG���',V�O���^�gQ��m�j��Y$4�[�4k-Ǥ�Aoݴ��q��C<V��EJ�t4T��ac��p��Ui?����D�,��Lz�0&�1�y����|X�&`�@�#nߙ��C�%߬�B �ǁ4����+-��V�}�G��c�vU+;k�C�n_�3^�Ю�_�>0)3�_֖�	FM��E��'˧�}4�Ŗ�)ly=���Vb��tN�M��]g��5�`�n��1����j�h�4KJ(TG�C�H~�n�p���)��	�.5Ӻ�o��������'��`=�)�Р'�RTJ��
�VYU`$�E�8Ҍ���C�3�J���Q�d��Q�5䝋�#,��H�,��s[e-�S6�4����Oof�(�����ִih������S��.�|P;�S�:��%�/_�9��e���h�dQu��h`>&� y�,êu�%����O}|s9x�O"ǒԈ�n�ǲ��@g��b��R�S_�UrB<q��Ѧ��s0$i�pa[��`�E.��Xol7z~\�,h�J���Z�L��9���X)ix����a��o.�{�����_Z)��C�
#��( 9$
4���j �fͭ8i���'ܱj�m��p�Ć������f�툇pm��>"� F�,�~PjE4�e�r�)n:�����U�4)�X�F�ݼ�P�D�.B^�[��k^��{��L�(1ٕ��Ðq����D)lXG��W�Z���x��O���W!���ߍ\i�ol��V�u���$�A�wp2*AP�XlxVHYEB    fa00    1da0����i�gg��"��ݽ�E�9�E��z�@�]Rx�x�D�?�Z3����K��:ԟy�X�fqX88�U��%�z���S�Ѯ��v�O߄	�	!����;��N+�׵��B��M^�P8�"q��n��F@Ҳ�� Vm�C������OI�ǐ��@4pa<��sS&��W�����l�e��S%ʠ+65���	��B|�R�_]� ����^ҵI?��d��K���d��GPfr�'VR!$5mrN���!&jx��l��/=�K{�Y(������Ģ������@ffj;���{-ס���)m�ec@d�s��q���
�9eAT_w���@^[!�&��
��3,��h�ĖUcģ/����yZ�FSn;��#q-��I����B'?X:q���v#*݃�Ip/Xs�&oxA�*Flح���ۂ�ɚ��B�vӫ>e:����E	�fՓ�1 �8���R��<&y���w7�<8خ��"�3���p��\����M����Ԟ�!4�*Cx���z7����Us�C����gB:^青�>i��+bvpUqP��Fy\T�hbY��Rr���,���(�_DeX��iBe�D�Me�T���# ����m?qy(1����n��
�����|��+n�	\,2��{�\����+�%���ī�A�́�ar�����V��=r����Z�۵��@�Ĩ�[�ѷ8�
){�$�gV� p�cy���+�ލ�����B��~��?��Vz�T>J��|�_F���F�O��E�Ov?* �dD`�>�2Hݣ�V�J���P��,�%W������^Uy9����>.��ʬ����d��#*ڞ#��C�����*�n\�g�����0=Er��D���}4l�FJ1[�|3#?FL�D2|w<.��mp1n��а�	���L'�����Lƞ,�3t3W7]�s�X7���#SK�� ��J�N'�6�V�X�-� Pg�)��Lp���m�WG2;�8�=��~׆���q��E_��V�x1����)������1oF����e@1�����\0�lm@=�IЙ��[#��|O�:ѡ�D�5�C�3���i>�<�8��+��sᰑ�61 �yy"'M�#@.�<p����v��S��W��M��?�4x\��TF�������g�:QW=����E̮��e��.f+�{�+��%�"��<�a�9"C����	��i��T	ly`4�:9�-~�
R♏��u��(1�uxT�>!��]ճ>����u�fK��<"�:t�ڶ�o�e�]���Z��o��츰��A����k�nV����P����4q�4K���#SD&��r���e�H�Y��1pO@���N��ղ�I�;�r�1�o|w�/��RR�Ş3v��qW�oP����]���<���[`��v��sʗ�@���y"aν�E,�K���΍p��jCV�H��	?o�����H�v�����������7+�~�6�}La���f�����U�ō-��'���)��j�U�}=Z�(����fS��6�y.1��	��#���09�s<��FAh�BƜ�>�[۱aZV�1���tV�F�o�������e���5*`aԈ�3~7��DK"<e8��5�|�,ڍu��k᧫Ts���R��J�1� m�Z<�g2��$v�2���������� ����E30�G^�G��Bԩ��6�U.>�{A���*�$3�A��(,Z��g���ǚ���.���ʲ�x|�QgK��qq��A�q��t9�����wG*�z߇�����.��{�û=�������5A��CX��r�h��P������ ��ܾ�]>:>���36<���~�^�@$~w���a� � ��V��c>H�&?3�K�.g��4��Rp���͔>'Γ�Si�f,j�y��g~}A9c��ɨ�Ek�F������C�H���		�Y��H��wdH�h�r{H[�P���َ��j.%���0N.F�_���)�Cj�4�\煆0�(�r#t2��q3~���ǲ�Y3�	��<�4�fe�_�$}.`��/�%�̛��mͿVpH���2����F	ю�gm~f\W�2#_$ɐ�+�	�`>���3���"ģ�%��93ϩa���d�E�Fmx�E����4r�A��H�w�D�&<�N�,4�#G�{�VHe�A�&㉫ D��AGULR��\�]�_���,����31���E���C)G���Y�o��sz����qЋ����n�d{| ��hŸ��┦��E���E�3Ɩ(D���:�������#0Մ���.��<�w�wQ�v(�tQ�p���n@Ie1@$BZ[|����L8��܋n,�Ϯ����P�%��P�f�d�
�`�8k�[Vݫt�=����KxEo[6
N�`��%��]R�&������ml��a�A&�no� (d�2X�̏Kڿ��h2�Bn��]GY5�t��r~�t�vx}�uŞt�լ�Ka�4�f�@dzE���0�9�ȓU��]'}\ӯ�v�PN�W��� ͙fԧ)����w���Wf16���:~��7�~	���2��i'ݒ�}�O���p�S� UC�;ߞW�hTf��]p^���D��b��2���)b�i�S���n~I'���W �ܖ�`Z�� j|.j�y�M���_0�\|I\�B�Z��-�X�cHK�_�8P��y@�,����#E���(�?�s�>��f�o����Z��[Ƈ�u���j� ��"usg����-��j�mP�	���;�G y�u��/�C��E<�Ω�_�����$9Dh��m'"E���L�ΰ>��+ۼʱSL�/X���p�Y"�B�)�O��3J���s� D�H[�gC�?H}V�����,�����:���`��/��T����ƴ�)��W�[��I�,.ڋ$� m�(Ѽ~ؐce��K?��@��b L��ȝ�4���.ژ��c�T���i�v;9����&�9zqĝ���&'�M��a��$X�-�a(F���!��2�*�����v��� �v�d32cfy�[/�̊�e[�;(���r�1��c�������Or����8
A?�(b&���*�-�>�o&�-�PT	;I ���!��%!�6� �UϚ{^���B�ᯊ����Ƥ1 ��X�}Mk���	���%�������\�שotG�5K����!���_+@����ҙ����dB�y"k=�*�)F ��I׉d�԰aJN����qE�{1*�zt�C��pnb]�@]2Q���	X'�H���'�L��pF�@��~7�	�����0c�� ��-MOdK7�(la�����6���4/�Y��
"����8�i���
���Գ�`%��!�����=n:��C!���&\}2� p��
PH_�~T<��T#*�O�/|$<Ǜ��U*�� ��M��8�}~���6J�,ԼV��Ue�.���$�k�}2zJ��SA���Z�g���In��BJ�Ɍ���n3m8�,�7�}��ab �su��k�4-5��G_��a�oN��YQg��������ߣ`�\��d&.>��.Ԍ-�6�Vh���.#nYM�ǉ�Ἥ��(��S~����{X��<LHGH.�C�������#��I\�l�q�'����p�<L�^�2g���K
Nq�seqB��	"���ݒH��.��<���;������Y����Ǵb��ծ��D��é]����i��$7'�֩n�7��_;�YJ��c/n{���ڒb���2����4I-s��-2���հ��+���i}D�e����^a�(��9�ض���zc\��sS��Q?�$W:Fⲯ�^�q���gq�
;[]��"Ξ;��8�p#RM�Sq�;��W=�}�w�%�	�J��9�4�t�p�B�8�T��@Ű?g�6���{��S���J��bKg�곞]�ˁV;��ֶMc�g�=�'�x4]��_�e��d׉I �q8�僱)��1[�9��i�B4��!c�|�?�����(���u�ȓWI�?l�d-M�*��O�zCR+�����BqyC�+%��N�@������m��:��L�-��.3�>��'��ޫa�	ξ����m�SSuIИ��cz��6l����Y�L/æ<�y�z��.HG`����We)ƞ�H[=g��YK7������OL��c��ÁfNR}�w�+��"�J;�@d��������4�Rv�XmF���o��@8a_�',�+3�O��^B9�@N�����5�w�D�lCU[�\�~h�bϚ�ol����2��W2��x;�
#:N=�<$T �H�P]��/�`v�'L�X卢�X��p���w����$�n�u�E:�}*�DNZqyXC���u����w��.�}ɽen:	&�7mI���j��+M�u��̥�%b�)�-��%UFu��gd�8�%�{���~�}��c��5����!*�?������N�Nn�vp�s�ȉ��?���2��g�W ��u�����N�%"u.��ݮ�ւs��l�bA�&��tc�]����÷�׈��Wc�����8�Mrk�bE�����'2ȓA�5�z㧟��Kp�<e�����Yϱ�GjcBu�NF�J�Lx-
���W�WQi��3�����[�T������v��><l5>c��aSn�QPd�ںc��	
d����Ԓ٤�ߏ����t X���Ys�\~S�:=PK�ӳ��KJ�	���r����`��~o������<訔#�{fo�ˋ�+��/#��	q�p����I�5!��BqQs?�9y3��h^��1���Ϣ6�<԰�tJ͓S(/5���I��M���	�<B+þd�w��[م^j��eVf�q��ZK"z[~�w�0��|	��틨������0�����+���g�?��K"t{�P#8bǏ��ELo-A����Mۂw�������_�߷��3K9���^�A�_J�y���w����ⷌhjH�JQ��W@�	�h����}�ݥ�p.(�x�]��8"�z_6#�т�~,G�p &�q�c7o��M�����.�1v*v��m���8���Q�vhCJ�H�0(��kU�cA>���,���[)�פ��ԇH�M�����E�[�ӎ��fn>=��PX����Sʓ�c��*�rR(|�����>�D�u�Bi�㥬�tR5��������Z�����א��XC@l"$�t;)�c���L	�g�����g�Ӂ��� �7g��R}�=�#��Gޱ�3�r?���N�134s����L��FK6�s
�n\,�+��g|~��ʹU��揸�V�7�N{a=����p<�랧ӆ��h���3�8/�~��ޅr���Z�	����W_42
� Oca;�YU5�qG~���$@�������bG�#���բJ\���V�*�Bn(P�`G5m��C`BX�|�fe9ڋ 3VE����׆�i�$��A!,���g�f�3�����ɦ?���N�_6��X<O���R(�١u"�l�i�p8<���iL��gJwE� ��ζ�Y���!;[���+�z!�e�n�ٖ[%���m0�uN�H�CN&�hFԉ�͋z��KL�(?v��D]l;Lc����&#ڪlN�3�9�8H���)�զf|ʏ�X�,{o/ř���tL��P��gÕK��E[��4V�U����X�X�m��&f���CN��H\�2���z���@"�
�����H�H���
�8��dؠ�B�)��T�a����QC�6�ȉE������/���#�bb��T��%��>�p��[�L֖��i��=��!���0]�����.��+/�0���uʉB#q���iv�ՙa�zDb�y�x�=�4��@�k�݇�-�Q��r=�ir�Qd�S|7{�!�'�쩭�H�ଫ�c�{S
��&YGߕ���T׾X����Κ�!)'�T:VC�e�&΅��}�[�m�m��q�!@b������mK�l�U]�������T�&^GAmߎ�'��6shR���N���7�y{�)��Z�k2��&��wf؀�r����%�/S�9Zs�h�˶���d��p���h[u�O����gxt�D��fz����澭Խ�E�1��QHI���9Od9���7ΰU�Χ���H��f����}�Hs'�ENӊW�Y�������s�SA�3Nۂ�e��/Zґ�5��ʴ>�fWO\@CK�&rS�!�f }tg/�}�J �㌶2,�t��2�|=Fw�I�w	��9:�{
�-&@�{����:TQh@��ˁ�8��4�^79�r��� �(v�!���a����c��,�`�Rpp�#�P�?p��D�+�Q_мp*Tl������f�O����.m�i`�P ���'�εj�U�$0����0���D�1VÍ��:S�T�p���sUE�Ha��~�K1�@9U�;��^���(!�������U��6Rӵ'e1�~.f�"�|����:����]�W��
(R(|sYqS�d� �my5���F��f	�uV�c�6BzyemO�VZd��D��ѕŤ.��Ğ'�q<�ům'�u ��r妡+I�Ldࠜ �xgT�ѹ�\g����XY�͔o�E����"�^d/�������$fT)kYy�O��N�$��ECX�
��SlG���>\���v5c+��H�F^�㘩J<f�y^�d�+g�~�'!�g�w�=	S��2�F�^%��{�b���n9��5S�	�f�e���}��o'�� ���c�/I�~�E�e�^�ʦ��X}��e(�h���>�Ƴ����[p�<���r�&6�?a�ցԿ|A�'�N�n�/Kf�%�@���������N��We��>�@��x���:c�'��ht�=8
��Z��}=T}ڝf����Lpю@WA�&a�����ͩ�`��s�~c+���Q�t����dV��T�F�D�Q����̾0�q�V�%�÷z4�"�H]�'�H��k-~��$+v̽��&-��E-�5*I`����j�@_���|~�{y�H}�il�!��}B�k%�]Y2�q����<D?�>o�ء�c�i5��?R��X�[���j��jEb�X���xL\�.��)"��MDV����7k�.���W�P7��wgM�CŸ��Q ���QS"pգ�.���%x�(ʒ#�Ex�[M�"��K� �3�L��6�)�SFK(�̛5�Q/�Ց)��"Q�YL��b;����Q�:��܎��>�؂V��Bn�E�GC�R�<V���09앪�i,S: ��(����\���~�Ʊ�j\��t;����/��d�K}��L���@��(#~R�w��M�[�-#�f�|�����]�a�yM��o��
2����Vd,�:����FLVU�����Bo�Q<cF�Ut�>N�"���#��1<��2XlxVHYEB    f314    1b50ݧZ�>�<�FAy;�o�N��x��>�)�,!%�Ho�D(a�Xʭ�eՌ�MZ0�:v])BE��Be�c��{&�ޏo�$/>J�F��>�vgoEg���&(� ���������{�1�i�^)| vk�Pg��WѬ�R�������L�3��B��Eg`C=���	.q�L��ߏ��M<jLh�)0�I��~�,��\�	�"Cq�%R7�@ϡ;�фs�,'�T }(c����M+kǁ\-���TD��:����@I��)��p���}������T6���j�k�oQ�6��F���~�]���CUV/⊴�{�I��s�L��w�;0f
�	��C�0�Y�VV��$�:ݸ~8�e]\SR��螢�&��5���aܠK6֬��D���"��N&��Ν�]���͔0Z�$4��;��iN���T��<�,�Y�f҇r���K�Lt�g�������]U��U�⿳�!P��ӯB�N;� �oޝP�ɂ�2�X�ᐜ�Z��k�`~H�Pu�<
�����<W�!U����Hq^-w�R�b����`�E�PE�H��S��ѥ'��BV����)�&����\��|��);?�u>&�����*���2jCX�G���.����U�V�/ou�R�;B%N�v�ɶ�l�W��� ίT�P4�i廤Z<��x-��e���p�9��FD�E�T�}�YW�FF�u�����2����u��z'T��Q�Ɇ~��Sj�z�G���7c'�o�L+���� /i
���I~:!r*F�N���+N��(G���c�G.]��y�����^�N ��zLY�!}���"N1ti��I�F'�\{$`=�^�C��9���m����ꙋ���zF��G���*(�Xv"�,z�݀V�_�%�6�+Q�Ճ��n����~y���������XJX3�׏�����j����c`C�����a+E�o�����IZ�}l��x^ˌ�Qm/PO�,�+W޿��Q#���0I�D�$�����,�~��WH�@�G�T�����;j��q���������%X�z����aϺ�d�~.c��=#U��+� X�a��&���,9��ʻ$���������l�fH<�Y�p���!Vm�b���)]�(L8�������V�kN������1��fؾ���K��c�LG�T�]T�p5J�tL��� +I���ffо�{��[�󷤕DϪ����Y� S1� ��Pѭp�E��%�e>9a���.��7:��UA��a��g�(l���بL������C5Z���0��B�B!�9�\�*��B�p��+f=�YЩp@����'�Ȫ~1�������p�`vPS�9�-��f�޻S ^�����?�p��M����dO[��s+_-���I����KK�c� �,w�,��`t��ʭ'b��X�E������`�=d����ޏ
?٫L|��qK#/�о��RڱL3����va�	|�� �i'
�ש�$�T����kDBcMU�N���4��UN����������=������in�ֳ���yP���҈�[����ϔ�>����qM*��JƄd�(:��i,�#�!^h��s�h	Ft��9�ג��N&����	�uQ���c� ������ 5��2I@��ʻL�Ud�(`@C�F�U&��e��Y��d"��"-D�#\2f3�-%�����a<H� �A5d��.��ն��ؕ][I�/��c�Q����Wa����3"f,8@II�g;�zv�)w�[�Xk
#�A����eO��Ijyp�]�\�$�C, /�-lN�/��d�l4M�)��9�tH�Z���R���\'k��h+C2<-ޤ�KIJ������j^�9Ԉ�2��u�r1?���5w��A3���;��0�:�NxϿs�Mf�k��L ڤ��U�}�c;?�>��c�E0R���n�֣%ڪ�7JU�U��E�=���:�n�D��`���� \U��c�|��~�D,�����)�xx��t�)��SB�,�^�~���L�=DX8���~�o/�Pk���!�'���&���� 3&��XyPu?N�@7���l.�����"𧐀;$��g�.\��O�omtH�*�%\�Q�ܲ~V��h n�	t]N�J)]ͮ��4�0Ƣ �1���U{-�z0�^��V�U�|f�
�)+�
1�"U���?�ڸ��-AԜ�L�6����2�Ǘs�H_��QZG[��o��0׋��?��\�}�\��X1 ���˒��@��luG�����^�"[��jH�4f�К�m��6p���T�Ö�?���?}��+��n7P�A*'q�����eepLFѤ��!��9PW��
�|bX1�ӆc��##N�6��t&��v�_u�9�V"��gDkvC����Ъ�ó��؉�:#�ı �,|�_���y�xCG�;�&�큰�;;��K��rF�LV������H�Z�T�OHᣐ��f�x��GyL�����ǂބjU��O^��Ү��C��:����8��9�.	jzF8�f*������CH��Վ�X���b2��к�k������PmYi�!���_ɇ��pX�'��/��p�����\����L�c���KF��P�h֍���;eOB}ro^��e�{�:"jE֙�T��7�AN�#[a"��ک�Y��K~��6��� H� Q�R�������jgU���a Hb��?�J�+q{���S�]t���7x��t~��!�)��Hr=��6S�1e������#�[,��6�S���>y���)�%�Ǐ���KT��З�d�Or�l@�g�
s:�U��-�����Z��Ƙy��f�����?ɭ R`�����펍�����ƞ":��_л�A����Fcϯ@ǗU�C. ��X��Y!�b�������j�T��rI�M�kԜM�G�c���mE����T6�5p:f�ҟ�߲Z0^A	ٲ�f�"�	-l�����y���{^W�#MAL���1'3���`d������5_YY��F)(*	e�e���g9�o�����;�$���I�.�L�%����	&�V\M���,�}9�Ǒdl�Vp�.z�<�M:��}џ;�iw�j}7)�G$sp��6ݙn{�*�P��USx2��T�+i�&�Q\T��BƎ왵lpּj
Flf�Qv�O4�A����inv�X�O����b���W�}40�~[��<�2�j� �)9����6���l�k:HQ)��a��8�e�� �X�J�(_�`}v�fTK����{j�L�b���_vN�$����y�m��h��H�� ��,^�T�N��m���:����y�W��u}�E5���3�I�/�Z��-=�m�~	2+Z�����4���c~��3�ו�|=J�u^;��_�m��y��,;ˇ�]�%=��:�2δNݵ�_J8M�S��ݡ}l�֔��|���d@{ZgI4V��[�ҩ��ר�K��,�@�X�0�8���z�6�%|�似va&2s6�s�$˜F6H^]�ED�959%C��H�9̶I!�^iQ�W*g��;=#am�=��H� �ǖ��k�nn���g���{���/֜�eJX�g��.���&���5 �(�Q��T�̷��bS5�b$IaE��U�۴�2��^����a���3�ѫ?V�j¶v@�m�gsw�ٴ�i��WE6�Jr�0;�cYQj��X!�����|U,[
�Nv�:J=�ᥡh����6��Ŵ����z��j�h�DEʉS���d�n���)�ֆ������$���곔�Ƴ��\X�r�����ԍ�w\x8��âk�`�X��_���'ʩӥ��QO�{���t�~�9��������^�|�=�	K�
l�rl�S�-��3?�x���9"d|Ř�a0����Gk# �+�y�SՄ{Mja�fs@is�Ɇ,�������5�?��ˉ�U���Q��?�J�.�F����}�.[
�L�֪ެ3s�D�����j����g��H_�d����!�����Vs��ͺ"[��� ��^e����.	T�ڥ[A\)m�T�q�wS_�:cÄ��W�۠�TBw�UL����&g�j��Aq�M��?��E?8V����~,�|)�:F���g�۹8�ڮ�	�}4j�W�]�%�t�@R89�ޙ0�[^XmJD˾�S���ˊǌ���ܕ�>�_��[U-Sh{���m�{��;؄�F��Q�O��AT<�o)�ϰt�e��C�)İ"�3�^��t4˿�aF[e��O��8�js��9�\��8����Ar]�^hc��4h��c�.>C}݀����<���8�k	Qn�R4a.#�g�}k�T$qM�l��p�*
κ75���tC��~�JS�4@(��wߘ���!��	d�1�8�Ë��A��E���:�f"���\�DX���7~s&iX�N�gL�F6���m��cU4Jo�.N(6� Y� !ۜO���l7��W[��j�c�b"�(ߑI�@���E,Q9�S�N�j@�H�hݗ$�[��"č$�.�=O��V^g���{��0��uz�|C�ˊP$J��&�`\f����ߗ`�粴����A�҈/�B!�����q&n��RQ8���]������lt!��Ċ-Q7��}b���wڬ�.-�A�C���a��ٴ�`!1�J��an^�궍p� ���(�����[�+�f�s���ğJ�3�0�'�z)�Dng�Ƕ8�d��������8�r�|�ꗿyN�Ϲf�J�'?eϝ������l�#�u{e�S����w�������u���!�IJc0]��A�u��Q���Mi�qc�S��n�s]�нI%��%��m)U�����&�ad�!p��K<��}L�2cܖ9h9�]�ץJ�9m,�k�y��$�7{�B�͓$��K4�wZ�f���1�4�~ge�7ׯt����/��u���r���������S�^W4z��+` �� \i]Y9-�x0�ߎI������\�d�XQ��oA�q����3Qz��V���t�NV�*�«��!��k���ǷN���0C<��At���6�]/r����M�[�րm��Z*�A�����Nt���6�/��/2䶵��K��z��c6��W�'u[�?��a��.��j�~4?De�SZ��<��h]`$�G�y�4�9iP��-*���q5��l~����m��돬���]&r����?<��^��&��c�������=�1j**Jg���Y�"#�z~_�%5��H�����NO�M�c>��Y�K.Qn��N���Ѓ(�Pbz9ĢR�#mS1r݉
�/�H�u�^�׻�e'ϋt�Bi�O��P����Pz�A�d�IG��)�|W�ҋ#�A+�~-�"Aj$����j������|���4~!xut�9�?5"�*0�W�m����ݢKбVO�(�	]�E ����q�*2(^�,ؽe�i�<���3�*��K�idG/{R��0��)	�$�) �G$�*�-V��7IΜ�e��ƙg5�r!���C�|M/+���L˜ٙ���F���2�_5M�Γ�+r�GB�P�wo�`F�Ç�$�#)VOO~�]S
Uc�m��������X�_v?��4�j?��k{��5�5B�h���Y��a( ���(T���`I���ÃVtL��5.M��~�Fb���U���@�fFh���Of��b�A�G��M�a��y&����\Mc�����T-
�-�S�vD��,*�Ƕ,�$���o��T�3-
��4��$�Ey���BL�>/�v �'��׻-RM��p������C�98�~J0r�zH�jd6��%]Xуf�����s������H���y����Y�Kq��zY�{����X\9�������:O��xj[�w�1���j��|�!��w,�C��0f����Ÿ���2s.���Z��˷K�?�<�E�6�IL���� h���g�9iٟ�v�&q��h.ڏ���)�q�������5׉)�晞웰-V;��uPb��^N�Yv�5�Ck��˦0L�α�/BL�%��¡L��ط~/��8��gW�G��y��bPk�g�LY��x0T{y4j^<��T�iZXڠ ���$�8��Z2�"k'��|�,�S`�iV<Ƴ�s�4�k�ѡg�0"��5)�s�462�v�I�}��³`�<��R���Z���0<B�u���������1Tv7�4��s7�\N;�tmh�63�[�#�{hH���9+;�U���´!0e+z�ũ+����?�hj�U�%���������ӷ�Z�Pl'�;��@$�2��?���W�Q��;�����O���b��Z��U���I3ZY��AԽG� [���b��t�G�n` ���� <�OP�M9���l$f�A�Fc+�%$t�ۉ4j�q��~�͚�*�����)���4�Ҹ�OiX��5A�%�@a�O���e���[+N˄�������b��Z��kBx�k�!p(�)�0{0���-z�K�E='U3#5��,�$����?\v����*^��hc'z�7�ؚ-�l�4�����������-a$������e�!��X4���J��M�x�$a`�f��>�ۜ���D(xW��'i]0�|��˶0�2wxN�+2jA1�g�Hg��?�h�tc�q�@l���͂�l�M��RG�r�g���.~q�D2@�^ӎA#��Qۈ/�
tC�B�۾����|�-xn9&O�A������Ҳ�2���'��l�[�M&�Y�y�$���g��t�K`ѿ+�ƙ�j�ɐ��ZnM�����f��yY���Q,ާ�*�G�m�b�@