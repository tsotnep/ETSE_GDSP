XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5��D��%[g�������jm�j��������ؔA=�%��i[:ϋ��ǣ�ܗ�����H�_!W���Y)��o��`!S	2H9��'�E7m�u��mL�pj���wy�g�
9ci��� T��_��hG@��'3��-;O���2C$�_=���fV����U=0�k��X$R"[�-Z^�Z�����ދ��Xw�M��:��W�,�VKH6��v��Q?��.��E�U�U�$쥅�����@n��l�!�}��L�3ބ���u�^Z;~�A�	����G��#[�6i)����ב�<8v!�_��v�8!	��r�E�=뛄��+7f����'�-��؋5_��JD�����I���Wȝ�� ��YN�n��Vl�\t @}�!�EO-އ�hv��׆�����`���[�+�N讬��N[�n2p���,�!��Η�!�����6#XV�j�׊SD,Qa*��3������l��ՀC�zQ�n5u��y>�õ��&J�1x0��ݶ�1n��-ԧг`�=z{I�֭���/ ~��D5-����8�����#�8aߙ����;#�g3kj��_?{�@�8bx՚Sq��W����cE�[�\����S*h�pYJx�T�2B�����7�igN��9�� տݳ�hv�u:'�ï7Y�j�/X�זD��:zϖ�ǵ	ܜ/�U���#XĖ�)m���]�}��[�e��Y�����pk�r��/a�H98����H�K��XlxVHYEB    9efe    1be0�L�� �_�Ǹ%��銽$Yׂ��.�F��C��o#�NJE#j�~��xO<�R4]�0;����9&����wi�A��J3ּH��{���"����AxwL�>��N<v�"B?�T�=(���f6��;���a�5�W���/gO���_&�h�8�ɛ�9~���iY!��m�[��v�\s�l����hyNX��������'H���8-��K��z 	��ɲ$���$\f�?��#M�ԐI��Q�[q�����j��]��J>�ӽjW�$N�J&�<�5���U��/�m�4�fP��K���QNG��F���`w�X���h���\	�~0�ʿ���2 ������i:��>g�&б���컹��}�������c��4"⳥MB�K��+��T�Ɍl't!^�
��j�������n����C #�»��٢<����ޝ:6���Mٶɑ�ｘQm�|�9a��{*{�ģ�v>��S�])�8���8�i+ =/tr:��w5?�.�E�1�8B=d�������S�\��2D۶���K��r�?M�zf����񻿒�(آ��,��8�97�'K2�fW����=n�"i��[��3�e�b��DF F@��#Z=�J���T:��1��D��2����Y�8��r�ʻ�P[�<R�Ϳ��V�2�n�A�w
4OD>��	�+#�f#��y>,D[��6���L	��Y��?!�bn���K����dظ��^�WZX�K���w�4!�l�6я�`�R�J:�iV�"�c�X�`�������`�>6�'�+���Z�G�������HI&�c%�U�u]���
�>�����7�e,�^�D�Tl�1X�ϱ���>��n��])���ǱL�|�*�Q�"	��ZFE7'5�� _�_s�PD�H[|/�r��Ιk-��{[�C�`+���_� �{�r誘� ]�zv%���OZ�v�K����� �`������kG��5��hv*+�4�Y���b�J)_���� �OW��@ފ�?����<P�C�� ����0�ES(��B�)�yG��/P�����߶���	��e3E�C�H����c~M�e��ev���Fy�'����
r�#�vK�o�����92B(�9P��	Ҝ��ެ������c��ϲA1Fe��h:A�d���A)��~�=o۾	n*��&|t��'�S�xw��'"*򝫤ꂹu3�=�)�֔�DA�˧2p�W���dkޛR���T���_`ݮ%�]�ޘ�斂@�R�Ye_F&�~�R���4V% ����O�U�[e�;���*�1�<e�$\粲�m�Ͷ$N��q��Ǳ��yP�4���ecw`��Q�hЍ��Mž`%dW���T��Md�4'!(T�Xͺ�P:���^�f���5��
{m��;�u/M~��]�]4fe�L!���Q8�m*=����
�]g�om�e�g�.0	.t�4$e'�%�bo��N��#�pQef��	��u�c㵣��~���IR1����� ����y�͙Fd���0Z����//��)��VZ� {��u�)�-�F�Q.3<��P�|�	�Xh�ۯ3���c�љd������8]hi�:h��N�l��5O7����C�BP��9�@^=q!;F-�_�BĀ��"S���/���D.Ee�d�<HGd���q�e14z�<���NU�7�~J1��($.�YJq��nq���v�깫Ұ=�I��3�^zş���9��h"��X�V>�nh����rV��o��;�X��|V�ۚT?����������[�<�3�rx��M���T��]�^W�ZƁS�Dh���,޸���h׀M8D,Jy�b=�r-�9G%�OƐ�I*9su&d�|�ќ(Ă��e�#��Ho'��iW�WW�&�	/9|�����)�F�J����#N"st�"v������O/��.nǋ��#���x�,��n�<f�!)������5��V�)��gÿ�]A)���7��'���?��[˝�J�	���3�]'�<�+�@NG�yo/i���.��4}�����^F�� iX�1���{�ѫ#B`i�h�c���#����q8�N'�/��2���,�Q	�i�ʦ�L��a2�P(�5�nW1�0fm
w��@X<�~=��?�P4�.��p��WT6�� �_@U;���q�]b�z$�0�U,e����&E9;7��K��@8�U�z�6��X���2<�)ޠw����+���^�� 4���9���a������@g���9(��k�S�	�o�م��knOј�q@t��`nN����n,��9XPo�(u����4p���������[�i�o� �h���ua��_~�>�ۣ���}�b�7��C�� �.`>���()����LP�A�OM�/��(����⁡UeC�UiBZ"s#�����q��7���yÜ�9�h��1�g9I��5_D�� m�Hō�w�6����u�F	���S9أ��%���B��B��Z��)4"$d�o�s�+Of�����ѡ'\7���JW��ķw;7];��'�7g�eHd���|�n��V�c�}�gԊ��jJܔ�`�=�rVP�ids?4=�50�(t��q��_
����Z���d$�fy�$��D9���>Qr�6�i�Y�or�k�V��O��ж�����6�8�!���8�T$���'K�`(��A�}�A�G
���?iA���3��y���6@��r��@���!\�=а�$R�7�F��2�)>%u��`�� �a5�}jF�Hg"�Nl�R�B~0����U�9�D�zC�eׯ����-�*���#�b#��amУ�i�n�{|��l%|�u/�s�U�3t����|̯`&0x� �"�h��Y�i���!����h�m[%�ի��6�B��o�p��;U�%ȗ��)W�5=:�"��+�g׻3��z�9�	��&ȭj���
�g�b��H�h�Ho�S@@��������'_5������:�vK�[tFToo�E��ˣn��s�?��R�������G��E��E%���%�:t~���S٭K;�r|���RM�j�#0W�-UF�H(f�6����L�=}�6�{r����i�B +B�$��$:��Σh#�~���RQ~K2�ZsC��a�����r�m�	1b���[S���b�^7�HZ�7�mH����rZ	�e3���Yޛ( ����t2��f;��&|D�{rӾ�'	�ث*w� �񟎀�ђ`-�H���Q�l\:J��+�<sB�Ag|{��./������C�������~�����Be�J�F4RF�)��5�C���u�F)i䭷N���{:cp�̑D�C�l��*�`VKt�e�74s��D^Z��*S&f��Y(��1�G�|��(X�n��Mn��a˹��b��:�U3��Cs�ijs��Y#�rqzٖ�ߎ��?�&�,D�� p	�w?������A�Ϡ�]�6�5N�>����2>�F�$'�~���:W(?X��MF������n��DW�3~٥��٩�%^'��>d�N��)p�qL�[��n�z h|�M��:�C�v����T�'��7�L�b-S�7N��F�L� �v�i�q
Yˠ?F�8N ^!9ב�M� \z��*BOѳ K��J
닱d	�(HtWů$As�Ÿ�K.ɺ�D��M��񠻯��2I!�/��0~}%T����[��y���gQ6��N��� �(M����2�M�|�E�Y��a5%���|�+֩�G�r$�#�	�#�H��}U;�;7J�� ����	[v��	D^%�D�L��i���,0�WG��Zt��k�)4�����:V��D�\(q7��dB�@x楡P���W�/9R]�����i!�QJ�������6eG���&=��<itf��)�ʽb�U7����P�]Jx�WO���Gv�9������\䩗J)K@�̻��_�.����3V� ��Tm��A?಼g.�w�BY�uTq��7��{���K)Mmc�T�m,�ga�ڧ﫛��A������]����N��@�0$b5]< p9Z
�n�('�e��#9fr���������>�{�c�A�����`�tJ��	E���s�;b���QEP�/J�M���Q���}Q��[έ��^�� ���+S9CGp%����4����UW2��~ֵ�w�5ų?�ݐ.��fi%AV[�Q\++��&\���M
�w��K%V��	���M@��@�!�K��g�2j����G^=�5��-�wD|��]����v��@��8�{��o2�c���=�+��+�H��4f�V?9�Dm
�:!��I�.�^O�pO"`�A�j��ƞ5�#ًjm�]B����<�=�!�3bX��J#%�^�����[yj@(<�jR+�dS�5^h#HqWi����r�dn���ӻ�DU���K	Ap�N��J��!�+�l6�k����J���D�c��}�M����߷>[)"Rn$	QO�B��mP�?_�b��nJ��Q�5S}CС2�1�:DJ�at��}� �O�?[vg�8l�][��]�����Z�����ŋ�F��a͵T#�TP60g�>W�VdFG=��Vn��[�Qx0�e�r"�o0�L��s�{�-Y����D7ɑ4�>�c\��}�
*�6��<�������?!���`�Q�"փ�n!�+MY���XH��?��m숝���U��ԍ�i�②������+���f7��-V�r�,���Mr�  �2*���2�=�nU��#Ė�sF �l�VQɡ����<R��m�����)� ���_\o�E�0�}�oz�ʛ�i����Ɔ��M�����ʁ��\̓Q�;|~���!(mt�����\�a��f�V>�46J��EhSK�uLB|�\�qQW�?��+o���<��������HawR�� Udk'b��gSXF�8	̦�}e������p�Nиv�|�^��h�dWe�b0���&e�a�Uϼ+�+_y��>Bi s��t�ɖ�z2E�̔΍�+�a*��I�X��?�6�A.����u.�����3�v�}#�f�F���)8A?͉�Z����g�bnh˃�Se@>Y����г��&�moA�ܣg�0Y����
(�v�$~3���R�`ÄN����[/r0i&��!:��|6Z�+��u,V�qC D���e��@�N:(!��f�����x0� 
����ܡ��:��$�>�qJ�[�Y� ���i��ne�EH��[bOꋰ�;��,�A��{���iO�;8���q.���DB�&���O>��Xꫴ�{�h�x�U�E�����A��BE�+` I� vԣ{�&� Ok��p�Y�%=%k�a�s��'g'�2;hS��+-���^�l�iR�Yrc�}����׎�3}�I���ް6�l�Q��[,~���Ƃffa�d���T�(3"���S?�.A	��hqИ�r)��P��3��N�?���S�F���S�mV�]"�`�5����I_R��rV	�&
�=�Y�'��!�\����߾ڮM\7�:u�pc�.���+�@��̉�	~0�N�q@n��2��EݳL��Q$9�:�V������Ȳ%�Ц=銊֏1h�����O��{�Nσ̎x����Ңm3�Zj�q��y�F� �cZ��-Ҫ�!��c?Up&/��|��ێA�~���$mW��􍶓�w4�@����()��a��]Y��)
N�Dx�kO>)�p%`�+��
��19/G;U�6�W<��λ����V.I���W�K�~\>G0D��0a���j����<�J�kjL`�L�o?m9n����:���i3�����mR����ѥ ��UZG�>W��vf��-!590u]����*]��^ۍ�-x(.��/��d�$`b� �jI'���KS���9�<�)����j×;�|?�o�q�wT(L~�~Ns�VB��R1�R�:[��l�0�-1¨�jGF����_�T�\o�VA�B�YAۂF9(m{4�����rhV<C���)��9���"R�K���HAo�e��]�������d{2P ��]9�� #R�+_.��U����6�%�����Y{E�w���ؑ��y����-�m��8���=�uLf�c&�s�Yu^8^��ƚ=�	���-瓦���S�T����1i����yz<:�Z���2Y�y���$� e���r��/y$ʛ�]8~^�|-Nq�|
�E�"qy�u��6�J@8�`%���>N��ڶ(��-��f�������{� ��F�.[�k�nܯ�,�GE5���v��F<��0F��k���1�iRj:w4���>�mI�nrLW�_a��υ�B/127Z�y5�ӓO�]��;l��)�L�O�o�����q��U� ]h�!E�������R�z��I�#�`�q25FA��	?Bg�9c��ئ�<2�,�
��r�oU�$��^��oZpq�W��ŧ��� Q����h"x-]J��9���g��2��� �a�Dǘ>Fj�O�4ٖ����g�Ⱥ4�e� �e�|����a��	A�kd�b����Q�&�mzV�?~)�����I%�n�qRf��{�(���b���8ڦ�[�H�u� ,>_8�����`鬡:^�e�2[D.6 �l���/�@>�lE@�"&P	31ƹ<�q��v?�I���+&2WK�X��]Q�Y���Ү�@eI��b��O͸֮jıߨ�$��~�n(�Y�@𤋮A^/�����p��Fc�^��K�e���>�:j��eY���7���-� 3���ŻP�ү�O�2o��"g]n�l��,ς���A��	�e��Q�ݦ���e+�:*�r��XaLꢩq�ի�wЦ{@��ͷ��=�c^A�C�R��?���%%9�(�N;����Լ$��<{���Mm��H%���W��ud