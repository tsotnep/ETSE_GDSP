XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����v՘HC ۮiL� �l�n��;��:����,�`�1J@��C�r�P|�!�O]dg��	��=K�)�	�M@�?�G�Cӈ�+2퍹�fJk�.�?nE	i��mV�m�!{t��1"j�P\���u&o�-[r��{w���^�^��b�EЦ �ϖ�ѻ���g���$ �2�/$��'�,��'��jw��[���>�p��H���~�"�_�0�^��?�ބ�noC�?�s��C�� ߎz}�����Ď�p��;�H��V6�+��
�M�b"C��Aa���P�ʈ> ��Z�S�\3bjr�^����r�(�Rn���M#�.�����*9�Q���/o	wBǹ�2,��V�:8d�L5�왬�i�����Ul	,�XC��"V�כY����kx{Ψn�+6����<��T��[��X�K���B��hn榶�(���=s�&�����5+I���y�E���C/T㡊m���B�n�@�����id\���9�Z�_��ɜ���������*�zԽ���6~iIC�t��x:P��:����k�s,p��֬���F))����z8Mj:=	�T}�3���; ��9������R	�i���.�3s�3!����T�E�ת�N�o}`�}3��F��v��9��=J
��(����3<G]��#��nevm�t�Hd����[��{�'���z�XD����@��,���y=D�n,[终��U(���_�*����Tˉ[:R���3����$+sP�XlxVHYEB    fa00    2910��^T<Ǐ8	`�E�Z��&��&��b���#��X�<�e�ل��pr��р$�*��z�k�̻�:ǁ����[��'�����1�L���g��M�i�0����ࡴ4�8��h��LI�3���X��|����JY�t9�h���9�[Oa���6��w�U����S��uC�m�@Y��Ma��ʓ>�N�z'+�F�J���.�|��/F��5�p�WEG?���m6�$��%�zt@�DH-,�M8GS7�;Q�0�LAǠ��̵����>V�cS`]��)��Љ*�a���\}�ti�T(�خ�o"��H;����M�p1�#�C��p�a�Fy
�W�d��[����H[`̝&����)tα����p=W��pP�����7y�ІVU�
r�I�bЭ �)s�>�6
f����h�S�`b�!!�!%٥�L�of�昦ozs�;B�It״X�0%"��޹���Fy�����!���ξ�@nc�b_mY�	�V#��
��r){����!i*�1���ϖ�=[1��(*��o��io{AF
�Q0�J����OJ^�R���d<˺N6�DL@�k��Xn]� �,�-�X`6�Tn��a�)U���L�d�n��u8+s�WH��8�?D��	�ߪ�����'v�<mG�����$з�1�1��j�J��Hl�M��EL����BN�"п1�����P9|K-�'J	M���(�m�>�ǰ
0�0�t	�hf�����B�C�#C��)Z(�ח�����=v�R�f��_�# uG���vE+����8^l�q�t7����e����L~o�q����h<惶Ġ�,sj,g���![����w:��d�[�"�0 }�`�4u9�����ɥcnC�IU�=(�N���׿�� �����5����ðX.i�#D�A]$�>�_����+%H�0�����/eD93#��_$��f	�)��"��E*j�Z���%Q'��Ĉd�s�_`m�/kTa�i�����ւ!w�};s��2
_"����|���Ч��P��`nKM�{�EyiZ����={�q��	�kۯ2���!\[�6��4l�Q+����D*�#��t�4me�,�&w��ڻ$�Ԕ�x�bg1.��g&����}�\n��t������t�����Â-c�f��oU?�V�o/6�_�S�=����x�[��-�OmK���=!���Kru����ɥ��=�q��?��������a�S�oH$�w\g
��H�՜��Ē�r 3$�R.�Q��4wC�Jm��e����.�3�R�u��6��4e�D���[*rK�*�[��AD7�mG��/e鹱�� h�xB�O�1mМ�t�+�xpM9��$�&�Y�� ���tG՜׻E,\-�z��	+�)T&���D�lHr���,�5�Hd���)[M1��H�:~���#�D8CUf���#��= %����Î��:���ޞ��4J��,�@Y��-ݸꔜ��hf�aj�uN� ����9�b�BJ�#$m�C<���WD=E˺u�ˬW��6��R��DU���a4H����
����H�>JR��oH��$��L�X�sg�3����f26e�|W\��6������c�(��e�
Y��Z�Ю
@���8 �H�P�#otb�2��指p$��Wޓ�wYuX���� �L��V�dKvL�}����.�䣛�s]2��D��\��$#�\������E�nK�i�`nV��Ƌ�9}]C�� ��h�'3���� VO����"�����*apꃜ8�؎���F���۹|����������F������ae���Û�|��@�e���|��p����KY�̝�F�3p��N��yveI�l��D�k(>�Hס�F NyC�  �}ʏ�]n!U,�Q�=�\(�Z�Zl�1���������$H2�-D��*�<��Ǌ��u��mq>��y�t��ֺ����1��G]k@�h�q�>u<��H-J�S���?D:n����)B�r|I�l�l��5��_��H�� :a>�sA n�;�ّUG�]n�xʯ!\%�̍{�IxH*�q�mM��C����h��.����mۤ	v�a�H��GZE�C0��4�?��zH�p�	� ��䓆B(˰h��X/H�v%�ߚ2� ;O�VY���܀T�c*#z�ŀ��@.x��F�N��G�5�T��h4��&?E�Ͽ)C���d� #�7�&��u��sSU��� [�<PC,�j��oB^��"�ox�?�a����6aOR���\��sC�+9�	 �p��<��쇄t���4M�3�]�Q:����΢a8<�	�����܌��������X*����fI�R���%pżL'ǲ�T\�[6B_eײ��zꭿ���}��H��:�Յs���SP�)��c�KKu�<�\���H��ū��v?Nl�PN��}*��J�*�S/H��H�]��%z�r����1r?>����E$F�tN9�I�K����im�F��|�����Q�؈�j��F_�zD���6]]�OviG�(tcs�M���'��f�G��ܨSങo@�9�H��E���6g3#R��W�o�B�G���D�׊h�����x���L����3P�97�{���6�����c�)F�����H53�n��3�;��~�fb������ө~3Ej�~�^��ah�D[�+(��7Iz�.�����h����U�g��b�Z���,}�U�􎥹�&7I�QXv�L��j�k��ϕ��q���O��s�5m�xbh���d
�;����v9Pv-�b�rw@�����]0�	W��\�k���<���]�����#��.b���^��}6����(�E!�؟��9k!Ő������"ɉ�lֽ.Z���5�$d'x���X�Y�]DT�V��Uixnq��,J}�9<��xY��K������M��Ob��z��i�AA��#��q������u�=�=�����q��V�$E!چ3؜�,:���k,�P|aG'"�`�qk�95�6j͠��#4���X&δ�R���8k�x� 1L�ț���\0�<�+�,�e|�Љ)�'Ŕb��O@~�bʎv�e�c|���-�%B��`/���3�T-4Kn�q�
c5�.�T������~z eh�1�����[�
�`ҧ4bI$%��+�i�p ư�S�S����$}�R�wQ͡߷�3 �N�ψ��U8e~�c��,g�jmm�v��,�8�mtF`mɠ�l��M�lE�'w��O��J�0_�y����j�kn���:�I��(�\0�z?Eބc(/�L
����Bؠ;����"RQ�f������6lB:d�@^M��Ʌ� I�'�F�'����%��%�y�~N�`<�C�s�IO�y�`���"g���Qo��*������C9m:�� s�׈�~z�8<f��E3�{�2o/��z����߱Q�G��W�a����鎙�=�E;�pߴy,ˣ���^{�vsq�O>�1�\-�]Z�vz�6�7��q��ݿ]iQ���$�!��I�jU��f��AF�x;	�.����/�����{$=*��e`]��z ����؝�0#�M��B<�֭�Ը��*�g�y���f\D#���2��싛a�q�����Z��EC'�vG�s�b:�9+uA��Nsi�I)���[pŃ 7[̓�:[͸�5�V���PF����l���:]���q#0�g)S����mA���I}e�4j#��q�(0
'�]�8&�oo��1W�>�������ӄ�5x��T��<s?��� ]����lI�ܛ'#<s�щ��G!���RxbJ�aP7\��1�AҔ��z��;��
�>r��D?%���`�S��3�i�r?���)�x<�*�c~j�~'���΁̭�03���>ɘD�1�{��:r(��\9��~-n�,E�sC+ݚ^�>�6b�ߔr��'���0��nq�=_��,Ϋ�9��KV���π�+d7P|�8Q��o��fug���̲]�ꈮ�����}m�0���VX�|F�)i<�������s�y����|<<���'�I�c��3z~�� .\���"�7jh�+��׶�g%�@"��.
�.��t/h���2U�@�8~F��}�(��8�#��y����6e�D-�� �����{��ҽV������O1IXg`j�$*�[`�Շg�jM:�/2�usӺ�v2*�NKV�ce�ò�0��g���\S����2�8�m�jON�;�+
L	U����"
������>�r���G{������W}U��޵�lg&@��Y?A�r��\�Dy[�<���傐���c�ڧ��G�%�y�X��l�d�
��Ҷb\y�n�W�����ٝ\���8�,�D6H��r�3{���c��H���g�E2��ˏ}ڀ�Ɏ���A+rb�h?���D�:��4��n %{r���Ls��?R���$BHU"-�,�bc�� >��9;�u�^ǵJ�Da �ĕU�0����=��.��gr�e�:H�l�?�S�ޥ�h0�rǝs�U�]�bR�p�~�������U6�1ֺ|.%}����bjcA8�3�>��U"�	w�ʵ��pg&XxN��v�S��Mv#`���K,L�����z��D1��|��`19��[c������5�HN����E���=Jͬ�&�q�7����{���v|?m�����~�{H��y��蚎L���a�r���o۹)�g+����F/(��c�'ͬ����=I MQ��"���3������Dґ^��=g�@f���@f�Q�x�	��hl�q�r>�NS�R�/�C~d��ڴ)6pD�+�	�L����l���[�]�����jܲ����0ԇ5���͛�$�����WB~�Ö8Ò+��Q�Ta���|v9��uXw����EQ�,4�����pme"襚ER��=0���DS��j������D�k	"Cj*��Ӷs��	����u��R����O�_:tmoG�B�R��$��b(?��#\A=���)���r�u4G/ $�_)ܩ�Ք)��%j+@w	/��vU���������{�GR�JL&u�*OV�4�zMݕx�G��t�����\G�H>�hTZ�Q<ѠJ�՛�����9��9ő��߬�_�Frm@��(�����_�A(����kk�t�	^�jEjI����;)��F�&pMa��_
v�%���-F9������b��g���S�rI��l{��+�8q�Bݭ�Xt;�]���\��@1�h���F
��#��Ϯ0Z�nx?�5۪�O3q�y!�0_>nn����&���WB���ǽw��l�RJ�}U�%��~$���5��=7���FO���{�Y2�'^K&O�����k���˱r�I�Cʽ�ދ�
�fʛ�tZ$���S.-�����f�SQW��
S�ut� tҀ*E�4�`T�=j���M [g�s7�����~�o �uMȻ?�PN�*D��yd��Y+��t��#�y�9!{�"���~&�����_�QL��Q�i�n [(:w��o����l-k��[O�������� �!I��%WC6���"�Y��v�ԏ�ýa\��.����N��xy���F�Z�8�PZ4f���o�w�����yVB�:���*� ���s�7��PI}
�Q�U���Â}�j1r�M x?SKl�V�A��N�f=?z��T��PC�X��&�ȱ Smy1�M}��mnk���*�� �LH
3��!���u,�T����>�s�%Jk4�Dih��a��m�oUp���ZZX9+fqڤ�u��N��N��k��h�~ȥ �SӖ�ƋX��Mɇۡ+N��,���ly���a����Ab��9�-�
Oڅp_���1��K�$���[M�A^8G�ti��
7Ϗ����Q�i�g���I9��G�S�ч7q
��y,�.���k�4��"߳f(Q�N �IQ�)L�
�#���ǆ�o*I�V���?@_�Įк���$�FٞU�
� ��)-P7���J-�	 $����]uݱ�B�,��rɞ)�TS��=P�����T�W��VT�ܤ����H5u[+�����̪Hɲ;<�ڷȿ��'D6g���$܁"pe�=���k�m}T����5h}��o}2�8�@s��5��U�N�)���;���f�Ow�s�V_B�s ������mC]��dH���S\.�[���ҭ��ml��0u�H��U����ɬ�jʿ�./����G�/�m��ʵ���8������}J�(u�<�˟�fe�u��!_��D��Ԓ�D����	F3�� ����`��Ԗ�rXv��L�z���Em�;ɇ�,8\��ah���l9�eܖf����c�rc�ߴ��t3�l����k�!,�i�s�EW��!�e|�e��X���'ʀ�T=?�^�qP����Y�쳧V�~r������&�GN�a��)�D�
P�2�4}L����9��rF���CY��N�B��y�:��Tkh�z����SAN�4�Kn�j����G�B:��ò޵+��z�SN/�I_qnJ�~bU�LMg1-�y#��t� ���)����4�裝�yP��1��1}�̼vE���Ő>U%��3��_T�{�l�W �N\[�4���'dw�2ɚ:3��6UR2rH���g�)ş�_ R���k��	6,�;��>��a�pIܧJy��78w �q�曺��4Q��a����[��Q�8�+g���D7U��*�St���gT5���]��Q���B���b�P�+�E��=����S�V��>[�����ENmƥ��L�iW!���&^r�q���������{2�  ��ա�GU�;���JUx������IQ]�Z˄�jX1(��@�����u��W8�Qg#���;T��U~�	Wܽ\S�Ғui�e9\����_�	�~���������,�4��j��0���^x<3e��SW;�&�տ�c�+�45Zm+���0��y��`��5���V�y�K
�
�M�M��%m_L��[��ذ8?����^�b��?�sM d�i6�y	z�К\/�vi��/ˌ�*}Z��{�
��9���[撇Ld�۪*��[��J�Y�Z�����N�w��AP������ME����x�G&۝u�R�1-���ZΖ@ �w�PƲ�߯u�q���u�L�ۨ6��f	�\���eB�p� �_���2L_*�+���s��.:=�Ȱ�4�A�靪I����yE�_+����P��Tו������2T��� ~�U;C����x�_��o�� �ᏩF:���4�7�3�+������(��4t̙�г�n�"bT�N�=ƚ�tc�����EHB1ɶ�_�iQ����� T�N#�w�<��;K�QAmX�l�5
��f0�M�R�@W�
#�F��!ڡ����R�>@���A����:�-dj�#ET���q��M�o��[e�_�My���������|�f����;Q},A�&������7 P�w����L���Z����E~ˇkP_���2G�:F �(tl'ƞy� u��B�����s�T|ُ�3���8I�_R��`��O�0r�}���k�J_�:ٛ˚�1�Z���?��h�c�����(K�=܊>�&D�K��}+����F.̭�՚Z3e��k�$�Wג_ B, Dm��3�+�?n�s6s�[+���N��ג��]^ﯸw���Ͽ� {xf�m���z�S��+�/þ�(kj�}�g�
p�u
��1(��`y����_&��_o �����̩B�hI4�g0Ȼ��JHEp1����,�"�	�Q�m�؊#�kZKmEO�d�L���ּqj������}�	�X�EQ�
�x �� �!2�)��(�bm����|v�D�B�;P���6�dj�v��ެ-һV�����п�ג�X{�ek|�J��x�/8��-ʻ�y��~�-N�8��\'!|�O\҆����s�q������z8���Z��g����u%�
����Ǖ?���?�P�`k�Jue0����K�����w�e(��r��Ǟ{�,�[M⢪��,�S�G�%�Osn����r.=Uߎ�> E�N�d�n<�+j��|�][i��1֙K��������:##��X���%^{�M�zm��������� N��<մ���{]��o2̳N��c1�j�j;�c&C�òC!&�JS!�s�32'��M"x��Y-�q�b�0ao���H.R�0*����Z���F%Q���@H)�||��w�w�w��?�������,�ڻ�� ��+@�z1CpO~�;�FϹÌ���%c]�A�����A�I��W��t��%NS�W�qֱs�Dt�1�I�{G�kb�UW���3����	6��d;�ϸ��iA��z���b8���-q����LF���`�v�?x�,�Èv�����O�~f}*f��[t�cN�RB����^f��6i�^�O��I�]�쁸�c�wf���b��1� `76���il}���0@l��*���6&^��h�m��#�(#:��RQ�v��'K�E�e���k��w^�s��퐩��D=�nq��A�&��fX��7!X+��d��({r�v�)���n%����U��3?��e��[.}o�R�� �T�cN����_�Ibo�L8�M��)��g��~'���{��1z�~|o��U�>&wu�u�`��H!Cw�e>�iw���#]���(dM�V�^�١�D�IVN��6��u��{֯�����_,D�}j�iNjB:h��C��u���m������!	�bT��Ȇºq�zMl6��~��~<re��t��W�z�G�jN�l&=	��͖(��5�8��
i�wR7R �}O�l�����j���	�pH�1tG)OW�����!������6.V��uf�^���|��z ߶���v���q�!T�"�7i��Ȁ�i�C�ڻ��W�,:mZ�w����/�s�U<�'�9C�t%���$s���#���&�삟�!�����,��:���T��k�����aD>\���QVPjD��Ϳn�Ӵ+�q����m��$-B@M�{K��#��-=_m��e�=Or�9��N�I���3�,�+�Ri���ּ�p&Mѥ�e����x[��.Vz@8CE�|tĹ��z�ZJo2ƕ?c�DE�.��,�A�Q��3�q4�Z��J�t.�x�z�;��(2w�:y��V:��}r!SC���,�-����&�=��Μ�D��(+�)�oD�	P�|��)�\�p��]f+�1+��.���1�~�v���������N�^]��L��x]�G̋k㢑9u�"�x�~�V杼RRS�׭��p�ǔ�B�"�!��<�O�,ط�w����W7�yE�H�6�3q��o�|j�y_T����z�}�[��e�e<�W��{z��0��б�;x@h���i��2��Xs�����N���O����7�!VO���8��ߍQ���҈�Bs�ɘ���O�;Z����2��`�?�R�yF� �!-�M6\i���"m�8��C�`���WP���	�ma�2N;@2����)�z���L0��H��2��A�bA-2�U��h�*;8]O�c���c\E ��
�+r���16gź���\$���Á[}W��Ӿ�O'���ԩw��7U-ƈO��̡��.@�U����� ZX��&+�r��_%��Q�ʆB����-� y�sC����ȨS�cb����<�y�;!�������r����j�\1l� ��
�gCN9��k�x�y�V㹁ޓ_whw
��^X�`����`���|��R8�����h�؄
.�4�.1��~�c�f�Aw�1�}A�aS���A+���-d��w]���,w��4%���t�h�I��ݿ����F�du:"�i''�VӲ�#����v�O�I���GDOb�ћ�0��W�kA�G���V.Y�RE�^��t^Y�C(�Ae�(��o�Q%��n@:�:�_�������x���E$[Fi��l �e�[;���i�X t����	�
u�F�J�ĵ���P�:�{ѿ��cH�U.��8���K�|���C�ܛ�x㋈Wd�z����=Z%��,V􆨬d̺�i��&��+���n��o��e��'~D-i�!��u�j� �C�i��u\�~[W����CZҥ����K�W={�[3:�e�\��������s���~q�)T������cg�����7Ri}U5*j�XXlxVHYEB    6184     f80��1_����/J���{�����"@ҮIf]~�=�����}�DydUن��O��G�����Pbj��+�G%`� �ba��G}��C�b4K�� ����q����%��E2`o���dY
��3���s�7�h��B����� �-�|����f���s_2�ԉȣx*D+�IC#���[�:�u(٬����ma�J�G���M}��[��=$� 1c�3"��N���"8�T3Q5i��s��?*��A~O�3M�R*���vom��2��k$b��ע�Q,u�H��k������R�-�;�`m[0q�t�#7T�[�S��:M�ވΉH�߆a�Cn`��p��\W��-�/aq�m��n�UF�0���0�bH��WA�ճ�>�6�
�4�%���Hn�6��U`O/a͟�<��hI�@��>_r��A�H>W�Б�+?�'�BP�/�y�Bw�? ��˾h>\b��Տ�� P3ko�)9��Q�ɜö��I�/T�)bI�}t�:,g�q r[�x��-�����>��X��i��|�<��������<����|;�+���x�Cn��0��'c� ���BǭL�;�&���8�����Ӵ�5�R���;HA��Wͫ�j���a�.�d�{��xq#d�3W�s�0��xN����	0|yT] �T��[����N-�	��M�YRg{O`#��2���"�e�g됄MA�0u�s��n5�0C2�Tݿ���<��L{;d�o��YLƔ[�3����z--�ֵ53��K���zdv��Ki肐d@�	�Vj#B� �A�k��Wn��i�aͳ����j�����\):����������D"��� �(=��s6���;>���apN�W���?��4�X蠃��F���!ow� �i3B���? ��$ ذ�\���A��/�}���@���wVj5z"�7H��e[��S.r�@rˬ�sr��%�V�ڃ��ȩ���o^��s�)n��.�$�e#�Q�񎻻�j�߯p(�0��,uL�Nw���YC�Z����PDe!﻽�[m�gy��*����v�p�L�k��p@,�V�Qg�O��=�z�O��������_�p$�g����mdߥ�G�׬��DY��ˣ�f߄�Q#4L�D�Z��~'BU -Z���^E^TĲ�����f�]���)5*/���RzT5M�� ����o����":L��S@wnQo�tIi���`	��D)'%m3���6����ex�GD@�ޙq]0.*�+�%�SkIc�:�5hb���O�f�x����Ƒ+�fN��Q؍S}T����ыp0k�<��z��j5�B;5-��� _}Ggt?��d>b$�o>&`�+���	ڏ����#M3>�b	�T")/F�Vi�C�������y�s�E�AEI�bou�#CgR,Љ54��cCX�p�,�}�r^CI�b���R���)���d�"<�!�&��"86䬛yW��e�O��H�gڨbA���Xu�K�c�d��Zs�elU_��=�sT6����d��"����D�g�����nO��[�w��'�z�	�D߯I�)��g��p�ul��]�$S`LtD�*���ې�EP\�Y�@qv�>�L�YL�[D���<r\�,m���#h��&	]��c��
�T'���V�cQqv�b^,m�x�Q��g*ʈ|kr��i��N�����r*ϳ�#ݛ�0��t��9P���]�t��:S�D��s0o����Nb���R�a�NW�2B��7�3�k��ޛ�c�x�E�ΒI8k�:�~�k��'�
��}�����]��dSy��=Ka��\ӓ.��IG���5�?Iadv�ԢE��ˉs��-}�l,1"�.�7�_���ё��v>�R*K�aPؒD�EPt6΄�|v��鼹R�aG�{���m*gC�F���pt�Qb�~Q�I��p�S��<��Lд��!9�'�\\��!o��8I�Y	��=Y��Oo�KIJ�l�,ί��U���=m��B7PbD�?�Z*��\<.c�@"t:GV��o������m���J:L5T�޷��}�&ȧ<[t?�1Y%g`s\d��7E���E^c��̱$�c�G͕c
�Sn]�{>��&g���%���x�ZJ	����]��=����F)_�P��kJ���[
���\���΃�V#VtVXƺ��U�Q\�'l�KB�d'��;��%�@�B^>P�	�7���iaG���ئ��b�>��\'�P�e��� s
On��4��J��̜ !�����K��1"�q��;y�������3[�LM��:�lU�}!u,?��7�,�Tz��L}|�2�;\=���
w��om�{�V��?��ڮ���AX���k��i퓞m�ֵ?4)x<�w��$!�����Sx�AU��z���t��ޣ�/�^�c�k���62�)�H����~��@�D���*��5g����_��t�� � �ږ�����	��.�U�;`
#U�O}d-���6r�X$#}�S����r���uH_�'��6��LjB�.��a9tI��:��C�oT�fA�-șp�i����t�\D���;ir�Y�p7OM�LX(iw�ٷ�q���.�v����;eK`���e�)����D�7��ѣ����8)	���a6+�"#[���o ��.�_|w��t�	g۟��a���@�X
��gYQ���plo�f<��m1���\�I�N`��{Sm��@�V"Q�5Q�d�<�Ż����	Q����������F�>��Zt��� +'��T�5y� �oؔMR���P�bRNzN��lh^����c��e��vt��K��W�cdRǭI��c5�y�WJX��>[���I����������̯JWQ�^-(-+�d�?x���"�'���Tԡ%!,�����@|����L6���̽V@��ñ�z�>�Ǣ�(a�D�����Hd�� �I��ͅS�u5u��'Q/���4=�m�wM�����#*e�b�.%rkZ�*"8�7�V�t��j��O�bˡVy\���lv���ڨ�Ҭq�^�O;�����+�.T����T{�@>���BY/w|f�[����T���7 �K����e��/踎������8��X��~�Q��m�3�<������3��j�H����7��φ�x��me�s�y"����k�r��b�Wú3rb��c���:%�ʙ�0�wi��f���ml�aDk��(���0SI�_a�.\γ�I!��ޕyO��.kJ��XL�@	�o�W��Իgt�bOi�H�f�T"�R�y��hKMv�m7T?<�i�y���a� �-�R����"YD�A���|�93+�~{�F�����oSVi?'��Bͨ �yK��ݐ��s!��MIC^9H$�I�"��^�0�hb�TV�F�C[�I�J dҬ�;aS�����Ȏt:�M��p`dD ��l-&/Z�z#���ୄ$�|`̯��~�
��.�Q;Y�[�g���Bf�A��g��E'ze[t������<��D�MMsEt�Xs��rdU�K�I���T��w= �J�P5E�xh�o7�g�f��.��ޡ�S|F��)%�<�ԕ�h]{ʺS���0�;%`�;=,,�(�aq�W�`Զ`�c�\Y�
��Y0lQh/���]N��o)�����m'A|�����B*p肸[W(����H:������/T�5U� ����7���76�������v�������8��V���z'�D!_���@���n�]�H�W oo���@�l����>HRx�|�G#x���X�Vp?�]�l��䢡ӌ�B����8R�2?_=/ƒ�җNFg�8�1�Y6	U]�՜�퉒�@�'���'�ˈ�� �LI���>0��طP��˽���uh�!������|5