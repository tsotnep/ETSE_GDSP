XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2}�?�J�vv-�>n�<	D<��J�����;4�p��"
юt��񉌺C��a�5�Bɐ��4��~˸����-��NXR��bW/nx��=ƨm��;D��6lۜ\�hS�+B�֡>X�[8F�׈�?��J*�o���vn6��~bmn����d���nk �^�E�C,K�DA�]x���k1>B��/yKM��� �E4C��g*gW �˝�����gO�+���,/�4`-�Zcًp3"V��po���SCa�2�V�!.[�B �[�Q��U��)/93�,u�h�u0ڭpX���{m^G>��1��Ĵaj~;�/�m��{2�NC�Ԟ�X]R��y"�����,=B=�P�r�ǋ�Hټ��/@M��|Z_l=��/�>"�bXL��O'�Hz�A"��n��N��!?>}�Hҧ�T�Hr�N}�����8C���:��Nb�;z�s�S��5δ���%
a�%�����S�}f|���HL�Ae?n{k�����}�,}��bUw7f�{�x��s|:W,�YWK8��h�������z��p}G2�G^c_ �_	^"���q$��T�I���w>���+�����1��w�J	[�F&}I�?E��|�r ��M������9���h�� ��l��*��*t�򮴟�����Fmy��F�A�)�m��v5��ɝk9��N��E���n�$�Sǅ,�h��&1Bs�j�.0}OX�,sB�uT�@�t@Ǉ�9�	!z�o[_A��?e�?!A*�XlxVHYEB    2e55     b00բ5y����a�n&~���-�x�/��H���ۿ�<4��[�2���p�">�ڍO�ii=⥤�.�^�� �~����=xB�*bM��f��&�����/�Q�a���+�hK��+�.���q�K�k:{�=�Hۈ9w��ᶾ<;Y�22wЬ~Ob�em�s�ak|-����\�{����|S��b'�>�V����w��\�t��-JL/;Ϧ�Anͺ�Z%������Xf�Q�U���#6��|��b{]�qy���Jpԡ�L��Oz�Q3���x���R��gIFy���ܧ��?��F�'�s>�����b��`l�����@�̜e�2w���p_A�Y:=mA�'P2�.m���yrr�
��Ĭ���Ƌg\87�E)����4�`>�[b���G^5��UA(�dBk�c��#�������qť972��O9�`�J
m!���u������8Hx@�X�&f�����ax1l>���]��K3U_�N��0��	
Rc�Lb���qE26|�����_Ke��(��5���I��y"��ҷ��m������7ݡ�Kbb�=.�ϗ�׳�3����Ѹ���#����똬�?��Rݛ��GEl�����J<<��\[�Q�9�:����I�i凥�0M����*l8yq?YFg���#b���!�m>`�9}96�foua����O6�25dҕ�q.G8��q!:܏ߝ��w�܂�3�*$��9�3�"e���1M(���C��<U�Q����u���"N����6Uw�`5#���D�|�9�Y��;��z���sU��4ӧ{��Xm�p�ܕ�&-X��u�t"��LMm�F�j�e?N�;�Ѯ��CT9�BG|�M �w��C@T/���t��q�d�ZT���:�AO	u��7�_N�;#cY	�xY��zjm� �F\�9�ݿ��5໔��5�¹�i:N��/2�$�`^u���Fp���@+o!��(��	�uU%�O�K6In����^������]���~�#^�7O	��������ؖ�,�����^_x�}#2��u��'bo6�������۱��r�W����fwJJ�:���X��Gb!a�^8��,(�S�&�E4ܾMY�_�#&�PƾL����r�VjMM��B���s��fC���V�6��Ӟ-zR�~��u:ߪ�x��G�#�u��喜�c�ԨlN�
�Y�kab�2��y�n�+�e�#lE�]ui>�2�*I��/���?�u��W$�f� ���O��ݖ�"��i��/��޸��$�2�>)ۅ�Siu��X P>5�,Q-��
{Xj
	�Ǐ��ݥA D?6M`�'r��aR�N�,b������]y�����;�cv��z?�o^ƨh9���Vz��`����^���)
)B�Nf�tW��1�4�l�d�s�`���C �{�/w���_����B��������V<����RB��y��;]��jS�/R�&��/��-����1A�.5Io���
 �#�C@��ئ�E�]PZ'�����}EI�<
��t(3e�f 0�Nt�!���k���|�!�:ay�G��c�Ԝ�맰U�ю��êc��h��=U���K�u9]��鑤�^��@6���bF.�?�P'�x����ni�U�Z�^��u��1N�<>�� �!ś�j��LЌ�-�J���T��I�1�t8� C0�:��0(���Y���{Ll�Y�K#&D=�з�D	��o�a����"��H�oF&C��r�1gv|�,��l\q?�(+���q�0~7���}Tl�N��S���Ǥ��+Va������J�6ODe��ms ;&�\�t h��\��H�O��TG�?n���7�A �*������Kŭx���Ļ�<N��c%������6����O��D��> �&��=!�Ƨz�k��f˫P׮e�l�|�(�lc�c��a%|S*}��>��=~!�Lv�O[ mX�!ML�n���,S& ���MN����gP�t�KM��}P��)so�j���;" �������K����䊴�d��o*��d�[����[�ȁb�?V��i��5���M2��2S9,���હ�� ����Q�nUɟ?����Sv܁T^|��2�3e����x�N�m:`�h�:P�17x�)Zd;VT��^�?GC|Ơ���;�e�x}��;O��=���8ɇ�?���*���nK����Q}���T[�J�Һ� ty�$,3����ӊ���E��
|6�JĒ�^3�3ɡ���͢��$���N8-�XH@P�%=�e[qf�h3��Cߎ���C��/ה,2~4W��5����X}��A��|�o�d�08�Fȱ�j�4����f�'��9����!�R[�R�b-��z�:��L�3�!
,�.�%�$�i��*��ť�����<W��R���A�y�/CO��^��:��o�8LЎBs9@����NS�ј�h\��y��cso1�m+k�GOB���x��7�K	���Г��{��Ã~�/����6gɅ+K`L��EZ}�&+[El���3�Wlc	7��� ��[T�{I�� rV�@�0�?k��F�|ʳ��>+hF�Mi��$2�#��]6��9�YU82���nΊ���B�:�n"Zd�ՃMW���K�3�\^� ��O2KzwJB�/�è���C��]���g�7��^����ON}���Vkk��+b��ۮS}� T)l�]�Xo-o[���b/�*`U�