XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E�W��!Mhəg��@A�0�����ǥ[����b�Z���,|��C�"u������/ yǒ?w���8��oW�Fޘ���-�^��n��"'�f����E�m/U^2z$��6kRLi>5�O��D�jm1FWs�����w���h.ҋ��p�ߘ�;ܫ.V5:E�X�_k�Sza�k45�M 3zC<2�î�C�c�*��C�BA�Vܙ�@1i��'qƼ�?��R��y���;�b��&����n�|�آ��=+�%�'�P}�o^oEb:슏[Ԏd��;[��d���=�؂3퀚�!�P���͐��,`=��ebe�����%;*����'������[��Cօ ���]Ej%�|���g�rH���l-?���A���Vx<��6��Ș��D�9���E���=�bA��I�e*�[A{��Yo��6�z�����m(�z�]�Q=��tQϖm�z<�@
��9UN��-���zޏ�f!P�؀Tc	M�.>ٲ�M����R��Y3�_1�l�֮��wy0�q�h���Դ;���	oxX����F�ږ�e������g*�v2o&��ZU���*�2u�0N-���M�IO�NCG؉"�-��\MQc8QM�),�m���bS 2[�,B����Mc�r�Q������N�`��ղrY��}�h���y�<<���_�Y.�F�P���Z��[B!%=tJ#��)-��cM�˗��t7��4��I�<��5�7�8s-�B/=W�XlxVHYEB    fa00    2030�}�͍�Q��=e���O'����)z�إn���i.�AGn��&�?.���;7�Pl0A/̰CvgKP�����H}Ђ>?	r�����}�����笖RF�U��j�(�T-���g>�9ADϭ��Q?#R��TĀ�v����ڞ�|í�[���E�nZ�@-�:���$�c�_��[�f��]�#aݕ�A����/$K��[��+Ei�E�d8}�Q�����Kb�^�o���� �ddw�h3��J��ވ��	�,V�K���d=�_S4�j�Q�ֱ{�Kg]�|���8y뷽�TW7�g<5�������B�U,=��BaM�r�,��c�SOwb��p�������I���'+��Ǌ�N����FT�Bo:�H�_��r�]������RE��Fz�@I$�>MgY��9�oQ�!A&��_�+��M\VD��mG��R�FF��DN����a��^)��w�P�&�(�O�R�4��$�5y��Y�a*���n�\�س��rwx�9�Z�}����+��c��u�����40L]�����<�e�;�w�Y����^��v�������d�Sﯝ�w�ǌ���a>�̝.	1�h�_L+j%T�
����X��f�/����_qv2�S��&�@�<Z�;Q���/�i�)>I�ĉ��C�Oo5jU�.t���aڤ��p�k�D�qLD ��?�9�d=KĻښ���5�ke-u���m�8�o�Xς�R'�*!^�j���@�9H%]B���H{y���W��f�+��V,!�f7*�`)k��[�n���ŕ���(���0#�?��KyoR,Up}1�<z�O"d��l@�v��UƩ��j5 �@�ݧi�$~���:�#T>�IF���m���Yc��PP���tQ�j��~[B�����F�oa�W�FVi5_��U?A���D�Ș�J��y�4o���1._w��X��ж�0������,�V�4���IE�7�0�<��P>�K)���`q�� 1n� ��6�*�avO	���������Ю�#J���C���r����8Y̩7�ƀ�z�}!�������������������Θ����C�73;�����v���Vr�*@EĊ4Jj�Z��r7�T���BkK�`�9[EDF���I;��Ȋ�}����I=�B��:Y	�`	2�<��ذz�5��=�^�ٵ�³����	=:,[�O�|�a�eFdf��:S�x:��2��������-g��\-�YU���J��?��i{�tk��9<֚J�����5�"x�M�m��xB{�p~͎D�Gǘ�-�����3�N�Y�l�������`v���B
����pш�J���`Á{��~���~���>1�	So�����^=��Bu,���wC����1\f���GwZd������ bT�Wܫ��X������b�=X��&צj;Y}0�-V�;4r3��>�p�|���%kyk~i�BPm���5l�AM��3����p�P����A[�@�$4]��|�Z����Έ�E��)Tv��44y����X<�q�j��9#�M<o��d����H��8�â��?6�մ��	��>�SM��z,�F�$Ts�s��i�݇�e�G�er>rN��y~�tn'��@ \&:���!����� �e��}I����&V����>�9��z�������>!�Z�o�y�:@rO�N�eW�4t��+�,.j���P��.I-'^��+8��j����2�XP�Z�����e��5о�7B-9o�ƍ{�7�O��s}˨b�`�������U9��t+�L�3-�%�K횜{#��y���&i��)\�1׏��W�<7��Q����	>l�-I+	��8x��e%��*1����P{M�2q,t���/�r�+�ȵ��F�ó/$��#�mM��D�؝v��\����(&X��	��厾';��X� /�z)�OJ�N�r2�Ͳ�v!Af̖�0f_I
Z��g�̘' 6p{/A�5��pd���􍠆$����^��d�ȱ�PiDO���p�Q������#�bc]�<a�B���HzUW�S�N�����Dv|nL<����N��i����2���R�M���e���`c-k����XI�Y�V������)�i$)s��*S��� <�/�qLim�,�N��c��Y�DX|7
���`���mpLW��l7�o7��t.�ct�j�91o:�*Ҥ��>:�`��7����{�l��pa(Fa�+�����Z�ΐ�*�KF�p5'���S>���%��d'%÷��
��V{�P�
�C��JdS(���1!�w�X^J�_х����M��/��F�`8o���Pt�S*�����ͥ��!]�.�2���$ؾ{P|��MN�F�V��A�Ω:m$��0��5i�e5��A�N(�
-WN��ޙ��W'^9�I�ܥ��sG�ah���1�;+�3��%���0�P1VJ/��z�m�dtC������VmЏ������f;�Up�*LZ�?ſ0 x=��t܌��[.��y�l,'2.���T��\P��)�b�,Ut�!�W�$�V^��<29�-�����e�Nx�`TDy4�T��� �Sځ[|���G?��,��\(9��%BsZ�V�� ��z:M1"��vF�6��3r.��)f�M����t�7��R{E%��+0rz��*���^����:����| ���KyFϓ5t'����5r4%?�4�]��EB�.�Ǩ̞[$.��C}VyF��4�����O�KbO������_�#^��Õ�t'S��G�n0X��H�Knڮ�L������j���7>��dfx��upԜ�f���U7@ѳ�# ԠR�A�D���d�)�H�`���V�z���hώ�-���Sk�O�,��m�Jѻ�8C�@ӊǚϫ���mk���U��)�|�b�Z2B�=y�ͦ��b��%v�OB�e�(�j��Whі�Zq�;��L	W���a6�_6�Z�yYl$}K��yhF�����ci��o	��m=�q1�UV�bM�z{
�p���k" :%1:w˺15�����Ɏw=�O���HC��B���1��N쩉�X
�[�#7��	���Cz���]+�Ds&������g��t��ߕ8��ӊ�����e#t-iՊ���J����_Gk��z����"��AEM`Uŋ�{�(4��r/T�򹶯�b­��� m��5��l�a^�5Q_��=�f����H,gT$]�M�r0��$e,���JtC9(�V�=��i�j��<u�6Px� x�\o��B�9�AT�H}��S� >��6�3�xoeS��9 uT��*"�a)�Lk�>i�tp&!��`���<�5��� �ֈ��] M�l�(����%6��-�̺��K�ә&k�Y� �B�YH�
j&W`T��>$7����Цqa���/y���W�����	���!�h�g_�D�p�؊�3�F�W�)�(HK��FxY[�A6�x�:��<��\�)sd������Pl= �5m�ݮL� ����چ��G���l	d�]C؛�I�Nnb7n;{��,��}$�`�~"�:��ۂ���`d�mP
�VC��P\���+2������r3]L9B��K���f�1{����D�K��L�	+,�R���}���}�������_ �7��s�-��ذG)�ᕷXz�&��w��)�J:�1��?b� YbA@)#.�t�L��V���jNR�4wYe�+/�H�� {�IJ�i�]�h�@��T�^�ed��S�܆�N�F�i1�kQ�8��g3��)LtO��`�3d�5:8�b]��G�FGVW����۔N��=�t���_��IBy�k����F�-��#}����$8ur�T,��ϸ4��$�V�|�N����R;ǣ]>��*����,E��m��l1��y c����Nā����+vs�c��MX�g|���8Q�mR���j{�L�__t��8pu��x�'<�Y��=S��t��<� 4(@1�v${��&��c���H�]��_no�����b��� �]Ч�#�t��x��?�';x�>�����p���k7�ȯDb�Q�n� �v�O�ɞ��*<�O�*rm���r��7���?
�,��A;�i(��h��tӯ����q�0�AF�/l�������q�LQ1��@������T�M	J��J�1��h�ݑ\r\���׬p4�*�6�$I���C4�s�[��(�����C���T�쯞J�$+uf�(����˻A����� ��������<.�x�q��>iL��_d��wuQ8+�Te�_��K����K@0(�j
_6D,�_б`�����3#���FQl�E��	Q�?d�F��W��]/rRܧPt-����]��Ӥ۾D�.<�N�7��@��U?�8X*>��w!��?)̈́����G�{y�G��Z`���#��fӢ�:�8�z������"�s"�$�K��4#?q��}���!�<C0#�!���F��8��\�n�=�j��ɓ�GA��q#\טJDg*�6=��"#�%����N�@�1�IvJ�b�d�8�.�I
��^R�To6������&��K��/p�ntm�>ԫN���J�Qb��r�^Z����4��5Zf�NXx�Q����ڬ!�l)V�X'�v#Cld,t�`^�7Z�O%�;#`LS`�d��̓��7�Z�j�����6��8M���L�	�E֪8�S�*�Ekio�cQ����Ⳇ\�bs�C�+��m˛����+=S(�c ���MM"dɕTx�}�y��Ը"^nvD�%��!��=<�W�{�z�$���;el�u��']� �2���f6�E��\aS���ϝ+����Mt�\���vs�Q>�д��,ě�1�LWf���G���W�+�{����S�/���%����5��.��{Uqn{��F=l�WV]��u�ѕ�S��D�����/�g�va�YLkP�b���;�L�33�p��`YT0=z���~��YH����(۽͎�5~N�IU�^ q��H�8��]õ�����,:�X�g]���_�6���B��eQW�H�|�׀(&�-GB_܍V�T���%4_�=sq��X0���3ЎUeA'V8�i#[�d^����BO"�fK��՗R��f���5��@���ܲL����qⅎ��u@4C�XL�1��\�*T�����1�q�T҈Y|�'�M�s�NZVm���ͅߘ�/l�`�m(R���QԚ0��ݶ��]�Vn�^_+��_yT��(�S��H�6��a�:t�퀂1Lh�/F>�w�%��������S�CH��\7@�- LG<x�8��w`�/�ʂ^��|E����0$���`��4�|��o7��'`���+0�%��g��������H��h{\�O"�?����У����x����=]
<n�x*�>��:;����MR�:���Q�cu�)j!-�k�b �<��v~��4!��"�Q(s���x?�	�]�;2���N��G&�n������0[�z$�3�~5Z��[�^��\s��FC���u�l-�21�?(�
5L+]�D��>��sY�g[�N �o�;��|��<��8�,c��� ��RB�w#�{A��Kp�E3;R���ɡ��Z)X�P7>��0�^I��7���hϣ����j���g-���&�1ij+g!���э��`w�8벧��%SPKb+a��ۼt�8��7����Us3)V ��7�D'���|�qH��^MWAs'��r;����~e�D y����c��`�(H0Cz���}T��y���������d%��?F�]z�K5�R��[������ü��w����1_?f`E��x�8�qNG�=_��xA���edb�ɜ�7"k��3C���~�n��ư��p�@���ľ|]в����@s��kG;��Q�<`U����d�B9(I���c#��65:��*QU2�(��C�M��+'�m��ѝ�
�πDI�bXz�-�H��L�!8�B���������*�	�)��)Y���pĩ��j�g������|��HK
gү��TЬ�;K��vR����v,��=��j�Mq��S��(���|e���k�i�Ev�޳������*�� e��JA2�낀���Z�!�s{M�	�eG�7���B��`Y�E@�ճ�E��,J\~�evw��M�6Ûٵ�iI�3�ǀ�xp��}^/·���Y�K<�l��"Y�~����>�G���DT�kNػft�v��p<�W��OT��BJ�蕒���N7\����5<�]�C�=?��H�-���`��0b��n�D>��~�����^,�Y��0K?�����t��������|��g3PfsE��b=3z��s��^s��r�'��[��T�ŚȞe+�_U1,��JF�
1v��?^��d��[���n"���?���%@6L<��,��g� ü��ǋ���\mpf���JuI�<U��(��,��;������U��T���>�~���=_��bSP��N�Di�����4� .Z_���ڶ-�ٺ�DO���.x�kH���0ů=yf?��Ҟ�ܱ=���O��t&�zIo�7 �L6�=�K}���9 �G<�t|���;ÿ���T��+�f�mo8B|d�| y�#��n�
�p@vICnz��-����q��L&^�"�hS����w�|uJN_�phApc#�>9�8w���dͬIA���$��:�i�������<�>��oi�)�7p��^��j�"�Jq+9d���.��W����\�rE�	D��Ӵ�x`��/�̽�/Z�����r����Ym�����P�@���q=�+�&a�KI=���L���ˢ��8�"��q�����E�k�R��w˂�0�S`�h�s�E�K���~�E>����L∌�b!WD7��J��p%�ؿ�z*~5��S��,Y�QIF���vg۬����(QRe���W�%V�;3iR-{g�E����E�T�����΄ނu�y��/��7���3Ͳ}g�=��i���eq.��C.���lk�C(�N��u�$�[�j� ���5�����k��Ь�����O�[��ڈ����,�LPyq^X��s-�4=|Oŀ\iW$�M�����G�U0������vs�O�E�&����r�=1�	��Hnb�{y"�4��c魁B�%6y��\׎lו�ڤ����g'E����%7�Y�9���Y���{��w	�/��
>���(��,��oN�݇1�=V�jk9=0�R�%�ӑ���mQ;ϠKr�޺��K�A�,�I�Z���#�r��6j/P����"�T[ð��*~ٻ�p�Q�7�Oh�t��.�wq�1�Ar��뙯��/�h�A��t��UYN��-�LK�����4yI��b��SrQ��MY�Y��B�y�������iU�38�LK�B1o��Z
Z��������@g+��&h�Wh�2U��6���`ބ0�R�5����_h�E��o�0�	���j3�����:���p^�K d�*�����e��U��7�p�!��Ȝ��ߒ?���w\aº'4z����Du2�Og5e�.w�#xi���%���t,��
�B�I����7N��K`{�',1u|�K�Ò�<f�)���Nԁ6!��"�5��R_�$�$�b��B�@1�5u(����@��\�E�}�4���f3��2i�ʇdt��u�
(Wͅ�>Pς�q/q`,�O!�M!�,������9t�r��LX��F,\"��"�5���F�ވ�Oj�) ��wD�d(t�����l�]S9�נ{���̔�PF* rtүZ{ڼ�����)��3�	��ur�HK+臨����|V���-�C%�Xܼ(ÿ�q%�G����Ǵ�g�i)�F�=�ݶ*����_�����y��ﲉ�l���ҳLeJ�zV[�
0d�g�F\II�$���ttb������mNv��q4�T��x����Kl��.����ƙx��*�H��������1o�8)��ʞ�N-�ۮ{䫞�kݏ���7��O���r�j��[Ai	�)ն^�LsXlxVHYEB    9620     d70|:2��31�߄�m���9q�ܾ)F0u�5���*=�&�m�IcMXG�/pOoo6�ξ��W�ۼ��O��3n�`�z�E�5�}��}+ �q����E��	�g��@2+���"�S�("vB��m��r�仏�2�k��0���q�*!��.ȳ)}=���ު���zؘ��b�"�h�
;k_��g�x|/�f��$3Ĳ������RJ�BAOJh�
��=��A�DK��2$���u#YQ�
�0,W���*)�fq�ld��}���U���s����h�$A��t�#Ǩ-oB�V�|B���LF��֖D��i#Or���E�Kiޓ�$ a
p���_k�&��2�����r�3�%w�졽1 �Ą*�����j�;J<���p��oӊq �iflC\���Hj�:d��c���py�ە�t%���j�b�];�o���U���y�,>�&�(�$�u֑;���a}=�	��;<�;�
��G�����5!C�� D�1JRf��@!2f���]i�L>��?��1�>�xM�`�t;��7/e�Ԋ[z�0݁w�~��FH�:Ҽ��|���TH���ֶp��̚���Lz@Pt��ѭ���!����3����-U��9a6�1[e��9 +;�� f�O�=rqn֯�/����ns�ITh�����"ӊ+�~�����:f`/I/\����W�|����t�g+�K�&�FA�i���`��b.��Z�Jc�ڬ��y5jjr�'|JFѤPD�͆���(A@����'I��y8�M/+�(D%( 綈�B8���GQn�<>xzo�,@��$��_�=��<u�R=g�������H����t�r.��7�o�݉���1K7$�~����M�V\i��K�n	���J+�^1�sn����D�,2�n�3�5��/^�d5��pv����L.F���N㩫�czC,���]����8���_uI/������[}�C����sc��+U�a����*�Q(�8���
f���ҹё+�Ьt���ks�h�@$w��X~E����P�UdL����8��%'�O%��AޅNQ����tm �I�à�g�"IR����"�O@�/�0T?>%
=�vМVʟ���Vm��/��P�FY��x5��t��lx` ��q{F��0�r��%���J�<p,����,A)��t��MLv��if�2�,�r��/g%��&'jd���7��憊kԳ��b4 5ĽֳN$�$[W��:��8�$ݫ�1�'�YR`�c���l���,�+E�hDEQi�R
ԂM��0@��q%)��(�>���@Q�������
�>��s��\��������^:7�ό���t�rk�˽��[�ā������5�KS:Sy�y�s�p�a��z.׿����V�k��A�l��s%���`�B0��nE��_�.��`}�U�����[���{�Kz@�6�>]��n��lDc�˓[m�����[oy��B�� �[�]v$��=(����L�s�6�k�Q>�� ��W$�c\�����?{T�q�?"�0c�A��8Ol����z<,� 3Ad"v�J�-�[��ʋ����N�����a�
?�&��tf��P�	ʣ|l}��k���/��f��s���z��ڟ��&�	LP����'�
;��Ӛ��'5���o�l6���&�2���UP�t���������8^3����Vi`u��ԍ�ɰI�/Қ$&F�j�y��"^W�O�t֨���*Z&�#��f
S	�3$�����}�<�8���6n��t�>���$�E��P�Db���t��n׬.��Kx��+���cP�γB��t/������7ð��w�]�FY���f�{���%ܒ�:�Xٞ�;��	�}>bˌ���bD!S���Nĳ�H�ģ0� s��điZػ�lG��ځ�ٍW.%�
=��	?q�̚��x<�z�u��A������A�)B'(��1B�a��6�Yz&¿�)BR���)IM�]��Mz��F�cR����Y������?�8:X� ��~�I����)[\�?~ۖ�R�ۣ�t^��Qyu�H���!嘤PQ���DL]R��Dҙ�b���Ң*�- u��a]O���`Ec��]�}$����O��9�(�B���K�J�V��!A�KLa��n�^XL!0�y�ɡ�V��X;I�1>�18��O�
�e	���
_'���X��b��/ Giܰ>�2����PIึbTnޱ6��LD��B�/�/����r���΢�"Q\�wl��ie�ͪ9H�LYt��m;�F�zJ>�����������G�ըv3�АO|*k�Eh��_��J��V���\������i�菽�-4�C�R)��ƶw�<0"c�e!T���8�u	[���t��(;�:�+��cy�bxZ���3٦��k�%�������ښ���Dq�cğr�K҆�ǉ^�4\ۯ�A���؎ �4��me���|�N ZF�zj����fx��)鬵\����$���v��
�
�]}`���y��Hn�C�#	��h���zd��V^�(7?�b�[��b�ܓ�� �4�O;TKY�x�w��"�T�,0�RkAp.�^�9ba�.h�&xk.s�e@�a�w�	������-�'`ўl4���Q��y��Q����σVP=�W�-��g��j���GK͌D0���/�l�g��(�?LA�m4od�$�݌�9���$j�,	O��1�(������^,]7F�O07sz����B���Q�T�	��*_0�1��C�U9�N�n�$��~����_���e�<��9�ѯ�v^%�C�F�;8S�	��$���f�����F��Y_?COK�I��9�8S�I5Q+EJ`0��;��oZ̢?���R�t6�e�p�#:tZ �@�z�w�`5�����I/�2�~3���HmH� /H����ƅ��i4f,e�Y<q=����(�5�NiaP�4;{��*�#1���4�\ɚ+��q�C>��,v�&j�w���I�l4f5!'��4/Wc�l	e�`�9�"�SfQpӚ6�.��x��w���Ĳ�0�=��^f�4u�JZCK��|��=�Z�:����f�W4"u�]V1�lƼ���=@�Ē[!��{�x�J��)^깿?�q��p&:��|3�#��%��}���-=�����m�L&�җ���˘�@��
��l�����#=�M���
��c?0�r�?1�ޥ�SM�ˡ5PS�v�LyW��Ւj��	�Nlk��{��Ξ{)�AQ�3^O�)�7��/�|>o�����y�LC��=4�7v΋�ޅ��[G��"�P��н.�=�ny)�;8(Iޥ��k;��J���1��8�`��?����_3�.�r����;�l