XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W�	������ !�P|L'A����n��g���
��)T���d�`7�)�E�خcw=d����o/a&mnY�5-[��x�	�.��o7Am|���$��)�������n�a��~Q(�\#7�ȅ��d/R `#�;���ef:��`k��i�$`�x%��/�rQ� ��ʆ?��-���sf��X���U8���վ��vI�/UA,[��tk'����8\0^"4��G�RpL �~���*�_���*�R�؀���) z� �&r��^�um�CX50QgXa˃�m26��gp'\�VƳ>D���.�i7����ˮ=p���_�Z<��k���O'����|X�����1�\���*?�j6����P�j�?"_�P�F9��9(�+/9�H5-�+
>���E�~�	-mH#w�?�j�4��x�K�ȉ��V8�`AѾYzs�����O�s�E��ĻF��\D;|�]`8���m�җs���h�,Ek�1n���]�jed��$�t�#׈�v�*<e�MnG�=z��2o�4�Ϩ+���O$���k?�^��o2�O�U4j�O�8��Y��������=�$ʺ�1�L	�.��K���5lu9˸�7C��\�Mvѿ�>���d6�9"���<Mp��^�:��F+<�W���@�^"ȱ��W%�G2��t�� C�?�'	$����d���MQ�cճ�����{���@�l���fsPoa4��e�9������Ԏ���n[��C���h�����XlxVHYEB    33bd     c90+�������qA��cK37-�3u��2k���@�z98�t��|T�hG~�5� ���:�qK��F.	]���]��a ��rjX��j�A������X��$���@?j<B5`z39Wx��3	����43g{E?�s�=D�]�$oCT�C'�sYZ�͘>(�*�9*PO��w$�&�d�a|��+P#n��Q�/�o�q�V[r�zu�
~���ON�-ԡ^0*�3LsAI�'�x{�ޅ�6�TyA-ij/�E�@z��0?�i�tu��J�y�G��"S�e�UK:{Lhxq~2Q8R��uW�ǩޥ;[�0jv n�+j* �f��-�� 7xCЈMv�#1�� �z�_�h;_�0�8x���tOqni�ڑ�J��k^�M���f֚��Y��;�L��!�X����ep��L��G�iM�7����z+���G�]q��
8ME��U+N�o�-�P����t?}����$�ƫ�)j�l>P�S�{�rqi����=t�2z0����;Ǧ�R47�E�"�����"<`H��5�K��)9��n�e��Њ�F>i�Y��1������9�J��k��jH�LVr3;�\�~W%⹵���lGP���4�ƨ$0� /�B�'rP�V88�u)b�Ζ�%���x�h�Yb�1w&u	?0���P�VSL;3�)�%� ��P�0&�[P�P�#4�cl��|���OURa8Ǥ��	�ʋ�Ѩʭ�{IR�țO�1�/`vkÕ)�y��}O��Qҙ�@�`�[9h1\,�_6]F��Κ�P&�(�/A����M�\�,n��p�n�1�c\�q�Ds�F��o�-�(%���kKj=�z��=�а*�#������[�)$^ �o�ئ��qZ7��~��[���b<�������nF�^��q�qJ�'c�R��FV�Fה�bdG�T'Ƙ��>�h�7�7�|w6�f�56�'���Z�l׍ k�Ɍ���3��إ��q\�S��������T1?��,��CW��
���N\{�{��b,T-E�6ͯ|��~)��qc���`�;�	_�/�!�4��}ɹ�<��apk�W�`��E$9W�j�q�<�I���K�F�?��C�o��U���R�V��$W�^�k�U�[��T7
`��W{�uܳo������</<-��&ӹ�8����[�3Т��� i&���ju���3�I!�/�䛆of_<0�~�F�!�r���,�9u��@xF�[�!�����k~K⚃� ��;t��'ӗ���kEhuL[��R��8���ǽD�"5L���{dWeK�D(^�B]8v�2��!?!!f4L��U4":O� ��+�� ������J��3����sx�������8G;O���x ��K���X΋Ԍ��~ƚe��۠W�⩚Eo�������U0��*�y����7��	2�e���� c����+�=k�nT�ϣFIx���Ѷ�X8=��A�ņ�M��ڂ�G	"�֋e��'���h���J1��^�K��+(��[F!��HQ��p�!ݒ��w���$H=�R��?�<% 4�}`�>��o�_S�@���$9�#џ�a�.VpƮC4�,=7l��}Q�!�TO�7�N/	ȷ�P�����o!U�by��b���&�k�̱�3�y՗����>�f�S���=Ό{A}��t�F3Wl��z-���u�3d���5hq�7��	��v�z��Q>瞜��*8L�N�:2�r_��l
�B�̸�-��;\��2���A��D�&b��qq��F,`�j5��a{��=�͵_�N9ѯ\Y=!a�:�3�nO��@�6�4�F�=2}�п7Z K��m��I-t!AO9�Y1����Ty�}ㄫ��t�-�2^
n������W�P�8n�X�*�{��q��=��qzGTb�j���TFU��M��hP�$�����(�	\{��Hbb��� �ْ�DR s#'ag#��*��f.�y�*�h7��p�]��}�3��(glVO
PǍIhN���w	�Bxk��.t"<7��P�G�U����7�:��3�O�W&�~­����8m����?ܒ���\�����>v�����a�I��l���OX�L�סDm4�9�c3ʷL_1� h�6��!4�M�D��2l���
��	�(���}7���9R����ٍ��;�<"T�����	չ�@����D�N$ސ�2��q���1it�;EYW~��1,���,@�S�{Sf����x7Ϙ��b�{XMF��&s`߲�i�wW�0Up�v�k�f�x��Ί��ّH�>���Lj��#����ۤj@-VD��)G��Ԉ-8*��۪^�HC�6P��@}'�# 7h��o���=�\����>`��E�4*��ˑ�!�)g".g&��^;&@H�ۚ7Em7�(�V	�2�����(E (k�7��Tȑ�|�yE!�R�!�z�]/����[���(��q�3;�z�����	 ��(ؤ.$���Q0õ��*�ɉ{�0�Dh��N*�I��
����A-���9�D�%��E[��0qX˞�>̓?p��T�<�0K{�u|H�mE[l��{���oc���������g��j��������CF(z��U���c-2�Or�Eyd-,V�B�@I���%W(�m}��L�mDP��z��Ԛ�!Ų��	=��p��	1�v;�G�5��v��B���ӿ
��h��۱Ǥ1G,qs�^��&�m����9����j�ƺ=]d����2�@���,�����绐� �vg���v��� 9���""�����?˓���9�5�u(VKy��`�'E4zЪI^��R�Rm�G���y����ߜ��0c���o曧'��έ�����drs}��RY�dr�r%q�0��v�l�R"��\[�'Yk䝗&�`(�N��(&�� e����d!+ǫ|�p*�#��%'��$�=����+�M�Y�$����Lܞ�"]r���e�>����Ë�&6-��=����GVwwԉJ>�ٛ���� Ng?O�vI��m�����U�RUƿ���{��!�A(���F��*g{B��u�l 1leo��QS9��&�]��N��μ{Vy�a��{ �]�*Ԡ�頻��������_
@������	�I� �