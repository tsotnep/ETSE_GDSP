XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ZC�;9	��C��Jx_mo��X���,��[�����Q�.��3����?[�j=��kF�U���^T2�c��Y*�4	��p�H��إw�W*[ 3��n�#f�I܇��p=�R)�Ԩ�W������D\|ذ�P��9��.b�Y����' �� v)?i��'�=*e\�7����t�=���K#�����{�,s�W�M3�g1��" б�(�����>z�2��/��#L�ߟ�圿r�ly�C����3�8 ��S?�M �R�ű�sS6b*s%��y�C��.����������4�F���X�]�.��h�n��D��g/��[�ׄ���͏��1l����h[�z�r��O5���z5�SS�1j�`C����t�*�r��v�V�z+g��r�8i�31���S�cm�ڐ�?�swu��{!�����dU��qO����x!�.\.%�c�(O��YH�@����q©�~ec�V�7���f�U�5�?c�bv�+|}K����6�8��9�>(��b��"x:Q+}ׅ�]�1�m�j���;^�|���[�y�=hT�s�@��4���.�#�$�+�09m�"o :r�^�V{���@T69�n4ʟh(Hm�31�-}K����c^�5�@nu5��a��;i�cj��S5�S"��V�z,�4VJg� ��8P��wR9���j��3n�DjX~��..��jފ��xQ�&��R�����a��|��,�}w�ɹ���KC9X��W/����oG2�u�`_XlxVHYEB    fa00    2d60�i��\�}!r���"b%�; ��
�-��.�殫�	n���MW7�.Ո|�u	�����ʡ�|���dAS�����ÃL ev{7���\MA1�[D����y����o�]�7zs��?L���<#�\���	ԫHn�Ү��t}j=�r���L��#�i���g�:�s3��	��%z�H:e��h��8�P��k� ӭ��J�D�V�|`�F�t����K�!��ō&������;Q�Wk�@�q:��Wx�L=W��} k��8v�Jz;+Y������ ��%\٪���՘ˀ(}�;7�����!d�y�� 7B�+������n���a�~K5�dH�^��u
S#��ID
go_u�cp�]���5�0B+a>���q�?���઀�X��F���a��]�!��J'�lx� 4�p�GFsd�u���*E�djx����[�kP,��#���0�6�8m~���d�D��&��}���1/5(�9(J�Q�ǒt�k%Q5�������A���u-�i�Wh1[퉭:"�B%n�FD=��ձCGѥ�o��L�u6.V�z�7n�:�����m��Gw�����x����9`	q�R���dG͐���	�H�IՓ_;����;��K���t��]��ܰ@�1�gj��h|�Z����
��n�i�?��Ax�P�S��ȗ�6�['��9Ö-{V�#zR�s������ʉ+�$��3�-���MQ	IA���)2\�B3u�M�W途��AO̐��z�}�T�=� ;��h���Åu���+��O�<���{4`�4u�q���~����Dn�t��[��Xzvz��;�ZU,j�?�r������>�f��DN�����U�
��c���C��F��H�;�mH<�N�y|��Y3�"B@m)�;�<��׼�e��D�'9�ғ�������e��}c�i�ko����%Fo}���a;�5�Y/㓬���Es����|�V-�����%�ca�Le.N#[��{��e�D���H�cK���?j�h	������
t�-�%��;�k��S#A?y�r���$.��<q�2���%�����Y�@�OƄ�"(�E�a�R$/26��;VJ���y���PnM`���c�0��l�L�Rs�ݺ]�.����W��r��B{M@�	3+$1�F吅�jh{H A�^�����o��sA	�s��$�qw��e��>z���8m5�q�4
��lp�t��ޕ1���Z�`Q�R%�AH���5Ym��ļK�U���C�F�ɧ�P���ቯ��߬�Kb�$���A�N�.y=z���UJ�U|�����<w�"�1V�U�ĉ�=�[JY�%�̗
�9���"�i��q��*0�@4Sŭ�g���JK=fw�lxZ��Y���;�Z�����m����N3Y��e�GtA_�y�\��|tč����T)Դ�>�k���Y�\!��ߺV���!�H��)^�iR�[�;�V��,��Z7���P� �5s���]SE��]p�L9
dzwQ�_��4�@TDC[	���M��}��g|�0�Z��n 
������V��ظh/q]u�A�a���9ʰ�򃪓��m�q(b ��-����c���C䕕׸�)2��4�P�f	�-w⫨����Z�#����)���4ݏ����H����+�H�4�ӂ���|}���;�K-v������tb3��*��	��M��;<��o�T#�L�IL��SWp�xHM��ح�b�)�Jb��^&2�$�{�?nq�CK�ݰߛD��?S��~m�
1��9�;�o��˽���S�G��c!¢ȱ]���آ�gk֩�|Qi2B4U��
�L͙8��YF���	��失/�
.�o�>�Hrx_������A�\�����kk�j�i��K�cu����XK�;#���$����d?��6,�m[��*�8-�,<��%,�����qHy~Q���i�� �#W��A��<��	y��A�z/Es�g�v�Z�Nl�[�.�|P�^֠=~�.�!�X���(>I�sn����4\4,� |�
��9/����e�o� ���Z�!��W����͓�p����P����{���w[�u5}k��׽;ܑ���u��SƄ���6�0�r�� �T���5����J�D7D.�DӰX�K�L����u��$��H�imF7�/Ⱦ�c�8�lҁ&�� H�ӆ�܅��"V?�N�k���ͼs��ONu^E	������-}�&�'%N1�Ԧk�m��On�K�?���>��sN�1����Z�H�eK\��A��l-�"���\@>�Se��%^r�yϤm�=\�w��:*oBA��%����� $W�YP�@�=�tP��ƪK�O��̄AO�F}�h:G�AS���rsރp�gv5�`��"�=Mދ��'�Z�-isF*�!��dE�?�bH<�rAA��r���=�L�!��p����)>!~x�ư�L�Y7Ⱥ�M�dgo����M�� ���w�E�5��{�_��@�Bb��N�=�h�;EV��8-"����+C�Hϡ;�R?��Z�r��)�~/(�
�FriL b{Wj�Z�d/�-#�M�TpX�j���yǈ!�?{��q���8�Z�x`"W��i���8���ߋ3 J���`�+��C��}�~���g�P�Kg}z��c���-�bvB��$��Z���3 �pM�Ӣ�Q2�ke��P��e���Z�B�^\'��}E���"�Úow쳢�Q$%8�����z=2��B���Fz
�-��V�1�Q���Hi��Ǝi�4R�*O�M�a�C�lK�ʀ�HE�,\^��ICTӟ��;�Tl�>�hD���P"&�/�vW�aZ�9Hee�.�B��#o���l���yѠ+$ۆ�ot9Y����� �Jv����7k��o:�T��M磊�7[!m� �e�p�F5^�G��t��Ž�rϰ�	�^Cs��߬]s(Sd@L �|hda�(a�P��@Ϣ��I�Z\>�d�������2��
�{��%9���G��Y_��KFV��A�e���=!�i���:+� u�S/�tu�3����-��0�F��w۰���
�����3�6}�x�6H̐�*^rX��F���
��z��1�a��KG.[��=�:��7�N+`�NϠ�eMLP4X���̝��ߴ�ן�����k�X\�</,˜���_SPE���nc�����c��;�t��!�ٴպJ�J��՗�3׿.
+ֹ��tNt�3����s��?��5�5��o�P�X.l�I��� <D���k��ӅY�@�8��+»V��hy�H$��o��157��g'��}��?�y���to��'j� ܒ�\;�<$�6���w7��J`!�{^r���k��!���{C���!w�0�m5(4U�s@	1���}��P�J��L��?1S�����$nb���cT/��&6pX���Qo��d�XXo���{��z�����Ep��D�(1ݕuUo�Deh���VP;}jX]�- k4G�J �z ������,{#מ�x�u��6^�7�hQ/��KI�q�ju��B����}�Gcd����e����T}O�it%��M�)��?a�K�Z[f ��s�(Yi&������4k�!a�mi�/;QG�wڞ�}4�#��<"�h�t!���t��T�*�{��yPR��m.��z�O����~�	h�o�r#����
�������1|�
"�Gָͪ��B=��B�G���?T7E,��;�Cu��b��a���F�F��8�d�:^���^=	�����'����S6�o�$a��� 2R��0 �1朗v�&��D!9����Mo�K$���ù2�6��>�(@X��� ���~�;R帝��B��n�������������aM,��J�
���c���7 �[56���P̢�}
`���/bx���ٜ���x/���⬑�R@�oHnP�O��c<T���Ձ��cLU���r�(F-���즁*Ğ�è����َ]f�2
����'��~4n|��5��ɹ��k���}7iU/>�國����L@"�f�������JTk&�K���&��H���D��E�z�X�e�ݙ.:_���h|�\E���{E�ND�X[���6>@�ۑ%u�V$^��d�����_Eqю����"b�mbC�;���|�6Ʀ�j�X���wg�p[nm̟[l1ƚSB��!�C���*ێ�*W�sΈ�B�'	�L�@�D���FR^�&�<K��(
Ғ�^���Q����xn~ê�W��a_6�(�;�>F���4����7�6��+��{Ԃh�����V�a�����6�,������[�ܻ9���zwq���F�������F����cZ�ٱ�k{M	���@��Ez!\xZ�G��8FP��]�v�Q�[:���V�o��؂���(zFY����0��t?�?X]k�a�� � ���ldWNRg�F��
�é�~bD���qS7֣c;Kh�F�g��]�)2�P�)T��w�S�т�.M�Oм��,wy7-��_)9��〄�Yd���U��yG"Y�e��Y��*�/p���D����@^��"�D�@N�������!l�+��CQ�O�'s�>+�^'b]7��_��u.�Lկ�B�3���pb�����TK��.��E*R�V��*������u$(\巙X2���dy��= 4�/�e�I{Mh�ha�N?�'d�����ڤ��}w��#��~����L�4
<�o7��T2b7�DQ�6�q`2.ݴ��8��|->y�����l�X��ʠN�
�Џ��;���1X�H�?O>~Pٿ��+R����-ӡ�`�T���dg��d6F�~��,Y�N�&��Q�������O;
��EV7 �ˬh�0�	#��+���Y�Čð"U����g���U�,�A^m�V�H��/���X �D	"�0����&�gc�R�����r������{q)z��[q���r��\7ڱ`��t�����"d�Yֿ��$��Ə!�~����1Ze��6U�5&�Rǽ�v�ky)���O�X��1�@&ư�n�	��n;��6]#�v����#X��*M:�>�������Ƹ��� �����?�U�r���q�e�=�Ql�Ǡ`���1�¼�4��$��0���3g��51�U"�wO�v˫����b6�ty�%�.��Ne+=+^�z(nQ�����p�J	]�ѽ�pn�G���m����V�(������-:)�.�7"ϼ����H�G
R���K����eFq
�O�<���ZY.99`�1CHG�p���҃�U`DIt��4�/{�2P4c�Z�c�E����w��Q-I�PJ};EbLR�
ȳ䵞`�صO�f~}��Z<�%�_�$|	�`�+z������s)�a_��!�b/9{r�D���c�v�{Ȋ�����e����a���,8�Oj���}}���-����]��m",��q���<DC�>��������A+��L����m��h\�^Go�5ܝ��EK��,=6�2$�[ۿ+ϲ�9XJ|�z%x��]����Sw���6v��@.%{}��0��?*�pY�ӮK�D$��3�h����r4fDJ��0*���K�Lz�,���b� ��u�Z���
�kb���^�X$?�BL)F��bOγ	|�R�o�Dk7���q�\A~A��� ��IAO��k}�{p�^C�~{�>	 �"��M��g�(�:|���_.y8x���	���X�wuNWf$p�����I���n��.�54�M\�\(�A�!��B�u:���юoK�.����6�*L��e-�/�e]GQ�G�_���gM�������jB�n�Bh�|���=��E�t?Dl�ER�ӿ?��Z�|l�db���� ���+�`���t�;P�%�_��T�7n�z�r}@�ĺP�x��2?�����(�I�B�1���ܐ��#d{�9������h�.e��O�}Y�;=��Z��[�3�O�i�����Zt/tɪICSo��N�N�J<�-�h��`}Ƞ�t[5����d��?sǓ	|S�B�0�(��f��uiv���,�k��F�]QK��b�����3|&eX���tZ�&����+-]S$1���+��Q
��[��E�:�U���*U�s�"�Dt��Z$�w*��_B?c�+¢v�����ЏH���	���h�[!G�����	�Y����@A@�fFo {7�x�҆֞6�6�\��Zvj6��s7�%�^� ���o�D��4��Z��Sm�o@�t���1\�y�d\�:2��z��%(B�#��ȿ��G ��%&�=S0LJd���5�X�e�[~ޢ��a�IB��8�F���μ�dz�jP�,ٴ~��;,���.�=�H!7���p��}�W�|YU�?�ru�H��k��O�?�y1��<�R���~�N���}���	��M0��wj�+~_�(��4���;u&��V�h�4�-��5.`��-u�])a'���_��'��|�f�o�=n.�[�G��X1?4OVo�>����o�Y����߈37�7MP���J%[����MPF�/�����;e����w('o,��9�Bt:L����Sy������q�8<�Q�`g5�Ԩ3�p3�����H����������
�[�OZ�G�W��aI�\��:VB��9�?����	2� '�:�mv6aV�
N?��$��8��U�,���q�����ϵڗy\X%/Y�$���"?V�Q�o����آ�<�r$�H�H�s���A�8���?��B6]��|Y�:A�`TI��G��t��X��Q�Iۢ�@e�-�ԵDfQF�dD̸�[�?�&�s��e{�{��`Hc������"���HU�%~x�FM�D&��Ln�w����O˟�c⇘N��n��ݤ
���-�R��u���ϣ!!�V�������
u_ ��B��{B�(���짠�6�VvdSw�N<>�������	n�Ly���S���Cf����`�.l��'�d��Gh��g�[%5��3d����gE�5��U���P�/>j��0W�T�vFWVG��Udb=�\�+5�}C�:���]<��������{�6�W��2�qe��=.,��m%E�ꅎ�uih��f���Z�%f�e5 ��?
f̉,��Z��1G�_-f�8�#B+`�'�tgU3��ݶ�!�Q�	���D��N\fżgu��5�1��wS�=5j\�\'��=&&k���d��P�Y΀��׏,�>�ݻ�\&o��|s]qu��dћ(�h7Ѡ0SA�K6���Q�԰��`@u�\�ֵ��s�%�P��p�����2�$�����5�������D���[>�A�e�5�"�۪������1�׌���{5D�sx�=�L���;����'�[�b<>���p�Ҫ�����@vZ���y�5ޠ�*�ӵi��P,ܲH�T�y�R�:�=���I+�ə��Ԭ�lh�V#��g�5G$���L�<}��*����q\Pn:n}�d�5Bq\Ov-
�s�y��݇
�M�$�AQK�9	2����-�dk��hUb|�y\l�6���RtKhz�������؁��(s����/%�kJ��p*��>��Gx�\x��g?V�}���|'��
�J���jgtX���l���>ML�]�K�j������!d4a��pD��ɼAm��KY�p9ۙG��RT�h�u����F|e˩?���@ڹ�����L��x�A�"?��,�+h��uŐ>�����X8-C�+E/OHǻ��Q�{n�vsB�A�m���Iǉ����0##�Q��~���<�<�6OO�ZK��`���X���+8c�S/�~'BZ��K�=e���9S׎z�D�JS�����rd,<Wٍq~�{Ȧ{��$�,��Յ�sy,��k�����|X�w۵/X4�����^�W��.fQ�Q"4��e{V/�.^��>���.�=��mϽ��O�x�[�C[h�Е�,�f�)�4R�u��\7eq��m'X�?��J�@{M�^��N$�$$Q�)Y�.ȗ�l�N�=3γb�h?���l�$(S�Hu.�����R\��P��(gF�؊�\���{N4�`ؒW�9�f�]ηR��Gz��u��ֶ�Օ�F��YD'Y)��R������n'Qv��Z[�aJ�|�wt���B�f�����F!��il�v,Ir�l��~�F,�9~ ������I�m�fp� E�nk�a��%�t.]�6�d�^�N§<��0;�-���o���y8��D�m|���W��,��~�;j��}�n��`:�B6>�y?��B�G�	�(q
ߕO�?B�N���g|�1�O���JF�V0>���*o����7��*�iJ�P�a@���f�Yd;��-j�iM����!��:���ʂH�K�v�?KO��Sp8�>��e�j��i`�����KvJeO裏�����N�[1���߃�5�9}�Eh�~����A���?�O�@GYwi�%�?Ǘ���Ύ�t3_��w��l}
��:�w�'O��)�ۚ����=�y���3YRYJ��|a�징�0��Ck(W�>�_�&@>߰�s� P�I�h�7�y�3t����V����&���x\ ��(x�EULyN�쯠:��יV����!V�R|��@���%����Pɠ�\cI�����V��Ҝt�#�U�dp6���%���ζުp&�R-I�i�e
��K1`5��j)��qpV!���>W�q�x��1?�f7��|��bJb_���)V�b��Hz����+�n0�|�J~@�ڕ鹷8��Gb�h��Kmò�G��4-v�i�#!�`9&��dE��㷒N�I�r�|��
�|�z����Y|İ�6X\D��Ԙ����j���JR3c���[�L@��d�c�[g_>�I������ns~l����U�M���?[��1���K�cP��q�	�`��)��߂�i�b3)�)�x�u�����;J���˔�Q����/ӂjK���Dd1�E�9�v�9�Ֆ�'��Hy+� �kϠZ���ql�<�������A+���p� "��ҙ�s�K��_}��,��T`�lk�&�+z-dH�+i!�i^��HF���e�5�׸��ȑ�S�t��uA�*����9�J��<?������_+�#CAH풳�0.&�IZ�;�o���XRT�	���2{�\�q<Hpx���6��mu]P)���,��0��!��*̀Z��2� j��q�G��L~XX�m��3��_�|��<���ʼ�ţ�)U���]�}���b��Zz�;�E1���0��'�(sN������D�t�X���l��pW�:�1��n2JxIq_)�]\�K⹲i��M��{��V䤺��M��i�y�Tu֗�?���q�60:�cvM5+��q(�����l���ʗ���v�8%����A���O�V���~����m�a9�D�طՍ���{?�lJ6�(���q!s&�2�4o3R�X�L���8��6h��/a�Z!��e���)�6�0X�]>��+ �O�uB�Ц��	�"�f(�C���f���v���WM$v�|���`X�~�.5hX�9D�y��xl�Պ�N4f�O�x�����K����u�(�G�rG��r��i^�s��fM����%A�"{Y@Hi���N�`C�ǯ�W������/�<wo	�f������!��GciJ|̛�	��P%��6� 6v��1"�=*�m��ڱ��&~�V�8�-,�cW�Y����G�ۏ-z��1�6�!V�#��x�7�S_����4X*?�����^���i���VR��oJ��h"�]�uě,(o�,�aS�-n�)������[�ru� <\��A3��Zu��cI�{�R$�V�#�Hb�$Q�5i����U� ;��1R����RDJF?}��ģ:�m��CԠ4�l�Z�zm瓷*;y�;p���ߪ�E�&	 ���]Ɠ}\������G��'!��<�L藒4ɗ��Ӗ��ϫ)yn��������飤����q�/��6ڜ�re:<�N�$|�b2����؃����4Cꪪ�0��s�e��SQ��b��<��	FzI�e�	R^�pVӦq��iN���C�߱�S��qP�x�����G�|F9-i��]��D	2r�I m�����A�%�罫�Y�^T�@\��i�I�w�����N5=�����l�Teh�O�;�#�������9ա�}ӝ�5���G�?B���y� `b�y�Et�{�����ٲ��N���q­�	��R���i8�+�S	5u]
g�A\A}W�pO	����g�՜�`آ�h	pY4��b�-��KC���O\�V��r�3���P>���yů�ݢ��)��]M"���YTc|�l�F���9��k�ٵޛ �[�fw,#M�Xs,MN7�^,�G;��Z��	��MQf���O��7*��+5B�[�B�C��x���b.��E�~&�`:���F X��0q���Eu��w{n����y ܔ�'E%!k���b�݇d��T��0��/K��^M�;S�WX�ޒ�rD��j�Wl�@���SFZ��p��$B�CK/�����n}�|9^6ϋ9�5L���dG����¯�rh\�����V�7"z�Bm�yͰ���v^$�n�B�W��(�օ��Jc߄��?P�
�����5�S0�J WZ���u)m�WU����hSjaW��pU&qm�\Pƃ��|��;���5�赂	�vbY)*p��9/��x�$�
���,6E�mi�Y�wpk�	Z�W�Ge�'��=얩5��/Y�j4uUm�< ��ľL"���_�R=��}�B=_�4��h�K�w�jW�CL�0�O[�1�A�/7q�&�^ɃSx�#Je)?	�|�J�y7L��|	^5���g�R��kx��8��X-:�Z�ɪP� �k�0���܎��l��I������Ye�q�[�Y�z����#��Є�W��瑿>ۤ(�-��� ��^�Dov`Q=�7S�Ȁo9������?C��#MD6Df�N�����R��f���r�1$�&̵[)���m��xd�9$��?�X�*#��T�����~ ��Է
'0=�g!�#($'��C�D���s.f,67�`�o�m"�t�������]Ы%\�+J�P���ql�Z����燼g�N��O��3K���f^�{��G��������[M|P��SQ'p������}>�Nq��Ɂ:QMv]sKpG��&ACI1��H5e/l%���E}�/�+1�W�Q������E�K"�X~	���hi�s������3lE��P	���TȂ��P�*��� ��u5����?�~O$���e9e�B��ë[r�XlxVHYEB    5914     f20ع�e�L
���A��:a�P1��IŰ� �w�6B���&��^�n�<U�2�1$��i�I�؁۩�2B݀A렂���o�G�6��b��ț\Q���LZκ�Q�?�ڑ/0�.��F�yh�> �<{z��y!*2>�9L�̀:��D��Ϲs&�*+҈��`-$˚�'�
�BČ��]� �f����.<�	}"F�z�\l�#/����7��$�~ˎD�w�+����(+������g�H���6B����9Ԇk���vs�LD��޻1��K��!�B�=ߺ\����y\WvX�-6h�S[6::���$K�+:���As�|1'�&W���D�vL��s�:n�l<(��b%���u�ަRM<gh�B���[8b��غ;�\��n"c�['�u�Xy+{T֞+�n� 2!H-G�z��L��a��3&v�c��G�l޽)Δ�����/���%�{/~��f�	���s8�+���w���W�&����ᠭ���������\��6o	c X�<ڹW����ÿ�K}�h�|rti�6uy�5F�	�L0�j�Ù�E��ձ��H��Q�����ܫ���-�r'd�g�h��N��|4[r����Tm&�w��%�W��N&%�G0X�+*�xt_������='Z������aT�P��6
5�xW�)�������������r�k����p�3�D���G���.G�3���-h��m�BEH99�����R؜�O�v��0R"����lݵvS�ߒ!\��u7�$�XU�L=���F�оtt�'o����ʅ��������7��^��Za�Nٯ�܊@�]X���X?��|�N��tE��:���5��jӊ�&��h尷��/_m	��YN�qp�����=x�R�H��L�-�ee��ï�4*�O� ��&j��7S=6��+��
¯��/��n)I֙�v�K����G1����H$���uLnŁ����s��_�j�ԏ���(Pf�nlp��������sS�m�B��x��ڟleơ��M�Q�`����@u��fl��M�l~h�^�-�A��6�r�+��eI���-Pi�Jv�����RJu;�U�O�$�G�	|�����$O�.��Pٖ�L����8%ˤw�<�t5U�ݗ�������Õ��2�a��x~Cf�md�n��Gle4Ш�t�J��{;A��d�3��E�Ydۂ����	_G�J>w܀�Z.h"Z�utK�����D�Z�x��G�E�E�%y}w�����x���|n�����u`W�2E0�~�%�`��Wpr<�n]>Û����:
�fZw��p����%�*�2q�nF`��CO������!�D�>-����؉솦��d����D�ȩ^H+kR=m���t^�w�$��ԆO�񘁂�w�>�w������'w5_b�� �fx��T��ٍ��}`N��/� s�[����ru6�ad���G/�1�����	_.��? ��x���!��V�5�ot�(5�ۍƨ��A:�B�E��2d��7*q�2a������g���?����\��|��
D�`IF���[�� �{�H�'[��a����5]</�尭z�
�����-#�^�EG՝P���dŰE��pFyL�j%%f�ijԄ���\�����BDmm_�Ig��`�E�[ǳ���	�Z8 /��rpM��~�p��O}�8$/y{"��㥌��B	��H��&����rwDM��Rn�ց��q2�s��a�+�^X���䦼S��5��//��������u���s���VK:�jr%�Μۅ��X�DF7��w����}��+�,"�/����<¼�@p�+�dv�t}�K�� �sm|1G�oi��2�b�!���a0%0��l�>e����ѵn0I� �R&O���Yl�ra��Q��У���30�r��.�|�|ς����J�~и�4��,2�[�r�4t)��>'9�vb��]ֈ��'rT����R��j�Z������j��/��T}̎�nYa��[��v��w�j�`97�ju�k`h����r��ė)�ύ���z�{�@����<�V�]Q,1M�$�N1@�N`dOEu(Uu�����n.naOإ&���dP��%k��ڼ�����efq��C�(E�`�N�U81��~Ȓ]���I�}��@�S���z�����<����"���Jr�C9gd+$0)��˶æ�Ցze׺X�n[}�d,Y�lsv�8fp��M:)���57��ׅ��L��y���ӂ�B/���?��|?�р42�t[�$��ץ]�zB<���W�vZ�ga���!�<Jy�w>i�!#2Bk0b�8b;���y9��TCnX�=�z��
F:@��G�][��4Ly�D�l�v�>�Q���_��W���e�����j���� �����<�a� ����pK�G��C	�n!eZv���{z���#��
�-S��hl5�����zݫ%���a-����hN+�Rg#�)�h�c����!��� D�CW�+��߹E��g��e�Ŝ\�c�a�Ġ���&_\�+���enB�t��&���"����'ˣ����ʹf2�Y&���a�;h���M0h�4����Ѝjx�l0,�˭��%����XlZ���8T��k!=�O�?����K�yz�I��P��t���&\x�_���.Z&�+�K�B+�w�C����8�j�-[��I�;A"8`gXjR�>�]O��I�y�c؆��s�,�v�϶�j�b��]S���j��U��9;�8��R���>�*3;��{��ԓ_�\S��+���9�௔�4��}m��L�e�c�<�7�%Uj�(,�����8d���ݷ=0N'��e� �Yc�٥�ƽ�x���ߧ����j�ŖO`;�oYj�p�M��УF��w�j5�.`�zc�	YI�Wc��R��5��0�Ք�K�ʷ���@�>v��{Q쭗�E �Bt�����Pz�ɞv<�;�!K�:-=��C�Qf��#K]��x�8���N�9�Q���.<f� �@���G0�������t�P��M�ֆ(�dL_�8�ʓ�CMw#�#���\��\����GTQ�t�X
D���gy>m|߷~RA�Q���NB6�n\����-�4��%�K�L�NU�6�Y�/
*���6�]���4�LOV����'F���i+ğ�B�����2���&��*$+:�L�9�j4�@Y*<�,�89���a��&��ɮ֫j������$��	��h�v/6K .��콠�S�9�� ����|�$l���tʰ���y�z��>Mկ0-�/	g������6��J'����e��h���ο�YJ@^J������)M�&��x���%ϙ�T�m:C�{D�0�}]�N>_NU�#�O��t\:�q�_��v*�	ɒ���nGQ�*ѻ���~L�;m��!�L��X��rl�|�<ȯ��^�:����O�^V:D��3b)�vt�e��I��~3*�á��1;�d��z����{mB7�EV��6,y	�j�a�KQl�ZȬP��Z˓3��97[���]\�qS��ғ���V���W�6M�+��T�zs�s�Ɓ���2�r�ce�	�Ej��f ��7?u(���-��47A��B#ԯ����kݳ�//�R7.��*�p�����E�z��^�T[�{e�{Y��8�|D�Lo�M�g�>�(;�#��Y�����;�+�o�ƽ��3��65>�qݐ�Q����7?�l�@�nZ�U��
�L>�ei���9��9�/S��R��#]M�+~�z���c�l�����P<��